-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    S_CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(7 downto 0);
    RX_ACTIVITY_LOGGER_pipe_write_req : out  std_logic_vector(0 downto 0);
    RX_ACTIVITY_LOGGER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    RX_ACTIVITY_LOGGER_pipe_write_data : out  std_logic_vector(7 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_call_acks : in   std_logic_vector(0 downto 0);
    accessRegister_call_data : out  std_logic_vector(44 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_return_acks : in   std_logic_vector(0 downto 0);
    accessRegister_return_data : in   std_logic_vector(31 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
    accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
    accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(17 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(64 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(87 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(71 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_3116_start: Boolean;
  signal ReceiveEngineDaemon_CP_3116_symbol: Boolean;
  -- volatile/operator module components. 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_r_data : out  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueMisc_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueMisc_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueMisc_call_data : out  std_logic_vector(104 downto 0);
      accessQueueMisc_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueMisc_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueMisc_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueMisc_return_data : in   std_logic_vector(31 downto 0);
      accessQueueMisc_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(103 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(63 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_w_data : in  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(167 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      max_addr_offset : in  std_logic_vector(15 downto 0);
      rx_buffer_pointer : in  std_logic_vector(63 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(71 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(15 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(103 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(106 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rx_buffer_pointer : in  std_logic_vector(63 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(7 downto 0);
      S_NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(7 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_call_reqs : out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_call_acks : in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_return_reqs : out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_return_acks : in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_ok_flag_1805_delayed_1_0_1911_inst_req_1 : boolean;
  signal ADD_u32_u32_1896_inst_req_0 : boolean;
  signal W_status_1769_delayed_38_0_1857_inst_req_0 : boolean;
  signal call_stmt_1868_call_req_0 : boolean;
  signal W_status_1769_delayed_38_0_1857_inst_ack_0 : boolean;
  signal NOT_u1_u1_1875_inst_ack_1 : boolean;
  signal call_stmt_1868_call_ack_0 : boolean;
  signal W_ok_flag_1805_delayed_1_0_1911_inst_ack_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1870_inst_req_0 : boolean;
  signal MUX_1909_inst_req_1 : boolean;
  signal MUX_1909_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_ack_0 : boolean;
  signal call_stmt_1939_call_req_0 : boolean;
  signal W_status_1769_delayed_38_0_1857_inst_req_1 : boolean;
  signal call_stmt_1868_call_req_1 : boolean;
  signal call_stmt_1868_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_req_0 : boolean;
  signal W_status_1769_delayed_38_0_1857_inst_ack_1 : boolean;
  signal do_while_stmt_1825_branch_ack_0 : boolean;
  signal NOT_u1_u1_1885_inst_req_0 : boolean;
  signal call_stmt_1955_call_req_0 : boolean;
  signal ADD_u32_u32_1896_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_ack_0 : boolean;
  signal call_stmt_1955_call_ack_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1870_inst_ack_0 : boolean;
  signal NOT_u1_u1_1885_inst_ack_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1941_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_ack_1 : boolean;
  signal W_ok_flag_1805_delayed_1_0_1911_inst_req_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1957_inst_ack_0 : boolean;
  signal call_stmt_1939_call_ack_0 : boolean;
  signal W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_req_0 : boolean;
  signal W_ok_flag_1805_delayed_1_0_1911_inst_ack_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1957_inst_req_0 : boolean;
  signal NOT_u1_u1_1875_inst_req_1 : boolean;
  signal call_stmt_1939_call_ack_1 : boolean;
  signal W_init_flag_1793_delayed_42_0_1898_inst_ack_1 : boolean;
  signal W_init_flag_1793_delayed_42_0_1898_inst_req_1 : boolean;
  signal call_stmt_1955_call_req_1 : boolean;
  signal call_stmt_1939_call_req_1 : boolean;
  signal MUX_1909_inst_ack_0 : boolean;
  signal W_init_flag_1793_delayed_42_0_1898_inst_ack_0 : boolean;
  signal NOT_u1_u1_1875_inst_ack_0 : boolean;
  signal NOT_u1_u1_1875_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_ack_1 : boolean;
  signal W_init_flag_1793_delayed_42_0_1898_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_req_1 : boolean;
  signal call_stmt_1923_call_ack_1 : boolean;
  signal call_stmt_1923_call_req_1 : boolean;
  signal ADD_u32_u32_1896_inst_ack_1 : boolean;
  signal ADD_u32_u32_1896_inst_req_1 : boolean;
  signal call_stmt_1923_call_ack_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1870_inst_ack_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1870_inst_req_1 : boolean;
  signal call_stmt_1923_call_req_0 : boolean;
  signal NOT_u1_u1_1885_inst_ack_1 : boolean;
  signal MUX_1909_inst_req_0 : boolean;
  signal NOT_u1_u1_1885_inst_req_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1957_inst_ack_1 : boolean;
  signal call_stmt_1955_call_ack_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1941_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_req_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1941_inst_ack_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1957_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_req_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1941_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_ack_1 : boolean;
  signal if_stmt_1814_branch_req_0 : boolean;
  signal if_stmt_1814_branch_ack_1 : boolean;
  signal if_stmt_1814_branch_ack_0 : boolean;
  signal do_while_stmt_1825_branch_req_0 : boolean;
  signal phi_stmt_1827_req_0 : boolean;
  signal phi_stmt_1827_req_1 : boolean;
  signal phi_stmt_1827_ack_0 : boolean;
  signal call_stmt_1839_call_req_0 : boolean;
  signal call_stmt_1839_call_ack_0 : boolean;
  signal call_stmt_1839_call_req_1 : boolean;
  signal call_stmt_1839_call_ack_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1840_inst_req_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1840_inst_ack_0 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1840_inst_req_1 : boolean;
  signal WPIPE_RX_ACTIVITY_LOGGER_1840_inst_ack_1 : boolean;
  signal call_stmt_1852_call_req_0 : boolean;
  signal call_stmt_1852_call_ack_0 : boolean;
  signal call_stmt_1852_call_req_1 : boolean;
  signal call_stmt_1852_call_ack_1 : boolean;
  signal do_while_stmt_1825_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_3116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_3116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_3116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_3116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_3116: Block -- control-path 
    signal ReceiveEngineDaemon_CP_3116_elements: BooleanArray(120 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_3116_elements(0) <= ReceiveEngineDaemon_CP_3116_start;
    ReceiveEngineDaemon_CP_3116_symbol <= ReceiveEngineDaemon_CP_3116_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1811/$entry
      -- CP-element group 0: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_sample_start_
      -- CP-element group 0: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Sample/req
      -- 
    req_3129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_update_start_
      -- CP-element group 1: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Update/req
      -- 
    ack_3130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(1)); -- 
    req_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	120 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_1811/$exit
      -- CP-element group 2: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_update_completed_
      -- CP-element group 2: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1811/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_1812/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/branch_block_stmt_1812__entry__
      -- CP-element group 2: 	 branch_block_stmt_1812/merge_stmt_1813__entry__
      -- CP-element group 2: 	 branch_block_stmt_1812/merge_stmt_1813_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/merge_stmt_1813__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/merge_stmt_1813__entry___PhiReq/$exit
      -- 
    ack_3135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_1812/$exit
      -- CP-element group 3: 	 branch_block_stmt_1812/branch_block_stmt_1812__exit__
      -- 
    ReceiveEngineDaemon_CP_3116_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	119 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	120 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1812/do_while_stmt_1825__exit__
      -- CP-element group 4: 	 branch_block_stmt_1812/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_1812/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1812/disable_loopback_PhiReq/$exit
      -- 
    ReceiveEngineDaemon_CP_3116_elements(4) <= ReceiveEngineDaemon_CP_3116_elements(119);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	120 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	120 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1812/if_stmt_1814_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1812/if_stmt_1814_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1812/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1812/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1812/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1814_branch_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	120 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (8) 
      -- CP-element group 6: 	 branch_block_stmt_1812/if_stmt_1814__exit__
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824__entry__
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824__exit__
      -- CP-element group 6: 	 branch_block_stmt_1812/do_while_stmt_1825__entry__
      -- CP-element group 6: 	 branch_block_stmt_1812/if_stmt_1814_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1812/if_stmt_1814_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824/$entry
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824/$exit
      -- 
    else_choice_transition_3214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1814_branch_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1812/do_while_stmt_1825/$entry
      -- CP-element group 7: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825__entry__
      -- 
    ReceiveEngineDaemon_CP_3116_elements(7) <= ReceiveEngineDaemon_CP_3116_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	119 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825__exit__
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_back
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	117 
    -- CP-element group 10: 	118 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1812/do_while_stmt_1825/condition_done
      -- 
    ReceiveEngineDaemon_CP_3116_elements(10) <= ReceiveEngineDaemon_CP_3116_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	116 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_body_done
      -- 
    ReceiveEngineDaemon_CP_3116_elements(11) <= ReceiveEngineDaemon_CP_3116_elements(116);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	22 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/back_edge_to_loop_body
      -- 
    ReceiveEngineDaemon_CP_3116_elements(12) <= ReceiveEngineDaemon_CP_3116_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	24 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/first_time_through_loop_body
      -- 
    ReceiveEngineDaemon_CP_3116_elements(13) <= ReceiveEngineDaemon_CP_3116_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	112 
    -- CP-element group 14: 	35 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	19 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/loop_body_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	112 
    -- CP-element group 15: 	21 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/condition_evaluated
      -- 
    condition_evaluated_3233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(15), ack => do_while_stmt_1825_branch_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(112) & ReceiveEngineDaemon_CP_3116_elements(21);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_sample_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(18) & ReceiveEngineDaemon_CP_3116_elements(21);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	116 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(20), ack => ReceiveEngineDaemon_CP_3116_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_sample_start_
      -- 
    ReceiveEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(14) & ReceiveEngineDaemon_CP_3116_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	14 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	75 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/aggregated_phi_update_req
      -- CP-element group 19: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_update_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(14) & ReceiveEngineDaemon_CP_3116_elements(75);
      gj_ReceiveEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	116 
    -- CP-element group 20: 	17 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/aggregated_phi_sample_ack
      -- CP-element group 20: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_sample_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	73 
    -- CP-element group 21: 	15 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/aggregated_phi_update_ack
      -- CP-element group 21: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_update_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	12 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_loopback_trigger
      -- 
    ReceiveEngineDaemon_CP_3116_elements(22) <= ReceiveEngineDaemon_CP_3116_elements(12);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_loopback_sample_req_ps
      -- 
    phi_stmt_1827_loopback_sample_req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1827_loopback_sample_req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(23), ack => phi_stmt_1827_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	13 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_entry_trigger
      -- 
    ReceiveEngineDaemon_CP_3116_elements(24) <= ReceiveEngineDaemon_CP_3116_elements(13);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_entry_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_entry_sample_req_ps
      -- 
    phi_stmt_1827_entry_sample_req_3252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1827_entry_sample_req_3252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(25), ack => phi_stmt_1827_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_phi_mux_ack
      -- CP-element group 26: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/phi_stmt_1827_phi_mux_ack_ps
      -- 
    phi_stmt_1827_phi_mux_ack_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1827_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_sample_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_sample_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_update_start_
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_update_completed__ps
      -- 
    ReceiveEngineDaemon_CP_3116_elements(29) <= ReceiveEngineDaemon_CP_3116_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1830_update_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(28), ack => ReceiveEngineDaemon_CP_3116_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_sample_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_update_start_
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_update_completed__ps
      -- 
    ReceiveEngineDaemon_CP_3116_elements(33) <= ReceiveEngineDaemon_CP_3116_elements(34);
    -- CP-element group 34:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/type_cast_1832_update_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(34) is a control-delay.
    cp_element_34_delay: control_delay_element  generic map(name => " 34_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(32), ack => ReceiveEngineDaemon_CP_3116_elements(34), clk => clk, reset =>reset);
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	14 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	108 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Sample/crr
      -- 
    crr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(35), ack => call_stmt_1839_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(14) & ReceiveEngineDaemon_CP_3116_elements(37) & ReceiveEngineDaemon_CP_3116_elements(108);
      gj_ReceiveEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	63 
    -- CP-element group 36: 	44 
    -- CP-element group 36: 	47 
    -- CP-element group 36: 	67 
    -- CP-element group 36: 	51 
    -- CP-element group 36: 	91 
    -- CP-element group 36: 	103 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_update_start_
      -- CP-element group 36: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Update/ccr
      -- 
    ccr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(36), ack => call_stmt_1839_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(63) & ReceiveEngineDaemon_CP_3116_elements(44) & ReceiveEngineDaemon_CP_3116_elements(47) & ReceiveEngineDaemon_CP_3116_elements(67) & ReceiveEngineDaemon_CP_3116_elements(51) & ReceiveEngineDaemon_CP_3116_elements(91) & ReceiveEngineDaemon_CP_3116_elements(103);
      gj_ReceiveEngineDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Sample/cra
      -- 
    cra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1839_call_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	113 
    -- CP-element group 38: 	61 
    -- CP-element group 38: 	65 
    -- CP-element group 38: 	44 
    -- CP-element group 38: 	49 
    -- CP-element group 38: 	42 
    -- CP-element group 38: 	89 
    -- CP-element group 38: 	93 
    -- CP-element group 38: 	101 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_Update/cca
      -- CP-element group 38: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Sample/crr
      -- 
    cca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1839_call_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(38)); -- 
    crr_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(38), ack => call_stmt_1852_call_req_0); -- 
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	111 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Sample/req
      -- 
    req_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(39), ack => WPIPE_RX_ACTIVITY_LOGGER_1840_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(14) & ReceiveEngineDaemon_CP_3116_elements(111);
      gj_ReceiveEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Update/req
      -- 
    ack_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1840_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(40)); -- 
    req_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(40), ack => WPIPE_RX_ACTIVITY_LOGGER_1840_inst_req_1); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1840_Update/ack
      -- 
    ack_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1840_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(41)); -- 
    -- CP-element group 42:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	38 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	47 
    -- CP-element group 42: 	49 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/barrier_stmt_1843_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_sample_start_
      -- 
    req_3324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(42), ack => W_status_1769_delayed_38_0_1857_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(41);
      gj_ReceiveEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	55 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Update/ccr
      -- 
    ccr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(43), ack => call_stmt_1852_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(55);
      gj_ReceiveEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	38 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	36 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Sample/cra
      -- 
    cra_3311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1852_call_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	57 
    -- CP-element group 45: 	53 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1852_Update/cca
      -- 
    cca_3316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1852_call_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	55 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Update/req
      -- CP-element group 46: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_update_start_
      -- 
    req_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(46), ack => W_status_1769_delayed_38_0_1857_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(55);
      gj_ReceiveEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	42 
    -- CP-element group 47: successors 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	36 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Sample/ack
      -- CP-element group 47: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_sample_completed_
      -- 
    ack_3325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1769_delayed_38_0_1857_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(47)); -- 
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	57 
    -- CP-element group 48: 	53 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1859_update_completed_
      -- 
    ack_3330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1769_delayed_38_0_1857_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	38 
    -- CP-element group 49: 	42 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_sample_start_
      -- 
    req_3338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(49), ack => W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(42);
      gj_ReceiveEngineDaemon_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	55 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Update/req
      -- CP-element group 50: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Update/$entry
      -- 
    req_3343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(50), ack => W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(55);
      gj_ReceiveEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	36 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Sample/ack
      -- 
    ack_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	57 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1862_Update/$exit
      -- 
    ack_3344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	45 
    -- CP-element group 53: 	48 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Sample/crr
      -- CP-element group 53: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_sample_start_
      -- 
    crr_3352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(53), ack => call_stmt_1868_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(52) & ReceiveEngineDaemon_CP_3116_elements(45) & ReceiveEngineDaemon_CP_3116_elements(48);
      gj_ReceiveEngineDaemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	79 
    -- CP-element group 54: 	83 
    -- CP-element group 54: 	107 
    -- CP-element group 54: 	95 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Update/ccr
      -- CP-element group 54: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_update_start_
      -- 
    ccr_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(54), ack => call_stmt_1868_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(79) & ReceiveEngineDaemon_CP_3116_elements(83) & ReceiveEngineDaemon_CP_3116_elements(107) & ReceiveEngineDaemon_CP_3116_elements(95);
      gj_ReceiveEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	43 
    -- CP-element group 55: 	46 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Sample/cra
      -- CP-element group 55: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_sample_completed_
      -- 
    cra_3353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1868_call_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	81 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	93 
    -- CP-element group 56: 	105 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_Update/cca
      -- CP-element group 56: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1868_update_completed_
      -- 
    cca_3358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1868_call_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: 	52 
    -- CP-element group 57: 	45 
    -- CP-element group 57: 	48 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	81 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	73 
    -- CP-element group 57: 	65 
    -- CP-element group 57: 	69 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	77 
    -- CP-element group 57: 	89 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/barrier_stmt_1869_update_completed_
      -- 
    ReceiveEngineDaemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 3,2 => 3,3 => 3);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(56) & ReceiveEngineDaemon_CP_3116_elements(52) & ReceiveEngineDaemon_CP_3116_elements(45) & ReceiveEngineDaemon_CP_3116_elements(48);
      gj_ReceiveEngineDaemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	41 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Sample/$entry
      -- 
    req_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(58), ack => WPIPE_RX_ACTIVITY_LOGGER_1870_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(57) & ReceiveEngineDaemon_CP_3116_elements(41) & ReceiveEngineDaemon_CP_3116_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_update_start_
      -- CP-element group 59: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Update/req
      -- CP-element group 59: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Update/$entry
      -- 
    ack_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1870_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(59)); -- 
    req_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(59), ack => WPIPE_RX_ACTIVITY_LOGGER_1870_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	97 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1870_Update/$exit
      -- 
    ack_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1870_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	38 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_sample_start_
      -- 
    rr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(61), ack => NOT_u1_u1_1875_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(57);
      gj_ReceiveEngineDaemon_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	79 
    -- CP-element group 62: 	83 
    -- CP-element group 62: 	95 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_update_start_
      -- 
    cr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(62), ack => NOT_u1_u1_1875_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(79) & ReceiveEngineDaemon_CP_3116_elements(83) & ReceiveEngineDaemon_CP_3116_elements(95);
      gj_ReceiveEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	36 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_sample_completed_
      -- 
    ra_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1875_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	81 
    -- CP-element group 64: 	77 
    -- CP-element group 64: 	93 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1875_update_completed_
      -- 
    ca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1875_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	38 
    -- CP-element group 65: 	57 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Sample/rr
      -- 
    rr_3395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(65), ack => NOT_u1_u1_1885_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(57);
      gj_ReceiveEngineDaemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	107 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Update/cr
      -- 
    cr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(66), ack => NOT_u1_u1_1885_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(107);
      gj_ReceiveEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	36 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Sample/ra
      -- 
    ra_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1885_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	105 
    -- CP-element group 68: 	97 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/NOT_u1_u1_1885_Update/ca
      -- 
    ca_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1885_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	57 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	80 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_sample_start_
      -- 
    rr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(69), ack => ADD_u32_u32_1896_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(57) & ReceiveEngineDaemon_CP_3116_elements(80) & ReceiveEngineDaemon_CP_3116_elements(71);
      gj_ReceiveEngineDaemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	79 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Update/$entry
      -- 
    cr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(70), ack => ADD_u32_u32_1896_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(79);
      gj_ReceiveEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	78 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_sample_completed_
      -- 
    ra_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1896_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	77 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ADD_u32_u32_1896_Update/$exit
      -- 
    ca_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1896_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	57 
    -- CP-element group 73: 	21 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Sample/req
      -- CP-element group 73: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_sample_start_
      -- 
    req_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(73), ack => W_init_flag_1793_delayed_42_0_1898_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(57) & ReceiveEngineDaemon_CP_3116_elements(21);
      gj_ReceiveEngineDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	79 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Update/req
      -- CP-element group 74: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_update_start_
      -- 
    req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(74), ack => W_init_flag_1793_delayed_42_0_1898_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(79);
      gj_ReceiveEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	19 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Sample/ack
      -- CP-element group 75: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_sample_completed_
      -- 
    ack_3424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_init_flag_1793_delayed_42_0_1898_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Update/ack
      -- CP-element group 76: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1900_update_completed_
      -- 
    ack_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_init_flag_1793_delayed_42_0_1898_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	57 
    -- CP-element group 77: 	76 
    -- CP-element group 77: 	72 
    -- CP-element group 77: 	64 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	80 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_start/req
      -- 
    req_3437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(77), ack => MUX_1909_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(57) & ReceiveEngineDaemon_CP_3116_elements(76) & ReceiveEngineDaemon_CP_3116_elements(72) & ReceiveEngineDaemon_CP_3116_elements(64) & ReceiveEngineDaemon_CP_3116_elements(80);
      gj_ReceiveEngineDaemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	71 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	87 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_complete/req
      -- CP-element group 78: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_complete/$entry
      -- 
    req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(78), ack => MUX_1909_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(79) & ReceiveEngineDaemon_CP_3116_elements(71) & ReceiveEngineDaemon_CP_3116_elements(87);
      gj_ReceiveEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	70 
    -- CP-element group 79: 	74 
    -- CP-element group 79: 	62 
    -- CP-element group 79: 	54 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_start/ack
      -- 
    ack_3438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1909_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(79)); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80: 	97 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	69 
    -- CP-element group 80: 	77 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_complete/ack
      -- CP-element group 80: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/MUX_1909_complete/$exit
      -- 
    ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1909_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	57 
    -- CP-element group 81: 	56 
    -- CP-element group 81: 	64 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Sample/req
      -- 
    req_3451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(81), ack => W_ok_flag_1805_delayed_1_0_1911_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(57) & ReceiveEngineDaemon_CP_3116_elements(56) & ReceiveEngineDaemon_CP_3116_elements(64);
      gj_ReceiveEngineDaemon_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Update/req
      -- CP-element group 82: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Update/$entry
      -- 
    req_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(82), ack => W_ok_flag_1805_delayed_1_0_1911_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(87);
      gj_ReceiveEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	62 
    -- CP-element group 83: 	54 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Sample/ack
      -- 
    ack_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ok_flag_1805_delayed_1_0_1911_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	97 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Update/ack
      -- CP-element group 84: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1913_Update/$exit
      -- 
    ack_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ok_flag_1805_delayed_1_0_1911_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	113 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Sample/crr
      -- CP-element group 85: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Sample/$entry
      -- 
    crr_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(85), ack => call_stmt_1923_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(80) & ReceiveEngineDaemon_CP_3116_elements(113) & ReceiveEngineDaemon_CP_3116_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_update_start_
      -- CP-element group 86: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Update/ccr
      -- CP-element group 86: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Update/$entry
      -- 
    ccr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(86), ack => call_stmt_1923_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(88);
      gj_ReceiveEngineDaemon_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	82 
    -- CP-element group 87: 	78 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Sample/cra
      -- CP-element group 87: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Sample/$exit
      -- 
    cra_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1923_call_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(87)); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	114 
    -- CP-element group 88: 	97 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Update/cca
      -- CP-element group 88: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_Update/$exit
      -- 
    cca_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1923_call_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	38 
    -- CP-element group 89: 	57 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Sample/req
      -- CP-element group 89: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_sample_start_
      -- 
    req_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(89), ack => W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(57);
      gj_ReceiveEngineDaemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	95 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_update_start_
      -- CP-element group 90: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Update/req
      -- 
    req_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(90), ack => W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(95);
      gj_ReceiveEngineDaemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	36 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_sample_completed_
      -- 
    ack_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(91)); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	97 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1935_Update/$exit
      -- 
    ack_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	114 
    -- CP-element group 93: 	38 
    -- CP-element group 93: 	56 
    -- CP-element group 93: 	64 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Sample/crr
      -- CP-element group 93: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_sample_start_
      -- 
    crr_3493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(93), ack => call_stmt_1939_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 3,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(114) & ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(56) & ReceiveEngineDaemon_CP_3116_elements(64) & ReceiveEngineDaemon_CP_3116_elements(92);
      gj_ReceiveEngineDaemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Update/ccr
      -- CP-element group 94: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_update_start_
      -- 
    ccr_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(94), ack => call_stmt_1939_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(96);
      gj_ReceiveEngineDaemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	62 
    -- CP-element group 95: 	54 
    -- CP-element group 95: 	90 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Sample/cra
      -- CP-element group 95: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_sample_completed_
      -- 
    cra_3494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1939_call_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(95)); -- 
    -- CP-element group 96:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	115 
    -- CP-element group 96: 	97 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Update/cca
      -- CP-element group 96: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_Update/$exit
      -- 
    cca_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1939_call_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	80 
    -- CP-element group 97: 	68 
    -- CP-element group 97: 	60 
    -- CP-element group 97: 	84 
    -- CP-element group 97: 	88 
    -- CP-element group 97: 	92 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/barrier_stmt_1940_update_completed_
      -- 
    ReceiveEngineDaemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 3,5 => 1,6 => 3);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(80) & ReceiveEngineDaemon_CP_3116_elements(68) & ReceiveEngineDaemon_CP_3116_elements(60) & ReceiveEngineDaemon_CP_3116_elements(84) & ReceiveEngineDaemon_CP_3116_elements(88) & ReceiveEngineDaemon_CP_3116_elements(92) & ReceiveEngineDaemon_CP_3116_elements(96);
      gj_ReceiveEngineDaemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Sample/req
      -- 
    req_3508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(98), ack => WPIPE_RX_ACTIVITY_LOGGER_1941_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(97) & ReceiveEngineDaemon_CP_3116_elements(100);
      gj_ReceiveEngineDaemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_update_start_
      -- CP-element group 99: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Update/req
      -- CP-element group 99: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Sample/ack
      -- 
    ack_3509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1941_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(99)); -- 
    req_3513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(99), ack => WPIPE_RX_ACTIVITY_LOGGER_1941_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	109 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1941_Update/$exit
      -- 
    ack_3514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1941_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	38 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Sample/req
      -- CP-element group 101: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_sample_start_
      -- 
    req_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(101), ack => W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "ReceiveEngineDaemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(38) & ReceiveEngineDaemon_CP_3116_elements(97);
      gj_ReceiveEngineDaemon_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_update_start_
      -- 
    req_3527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(102), ack => W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "ReceiveEngineDaemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(107);
      gj_ReceiveEngineDaemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	36 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Sample/ack
      -- CP-element group 103: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_sample_completed_
      -- 
    ack_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	109 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/assign_stmt_1948_update_completed_
      -- 
    ack_3528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	115 
    -- CP-element group 105: 	56 
    -- CP-element group 105: 	68 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Sample/crr
      -- CP-element group 105: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Sample/$entry
      -- 
    crr_3536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(105), ack => call_stmt_1955_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 3,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "ReceiveEngineDaemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(115) & ReceiveEngineDaemon_CP_3116_elements(56) & ReceiveEngineDaemon_CP_3116_elements(68) & ReceiveEngineDaemon_CP_3116_elements(104);
      gj_ReceiveEngineDaemon_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Update/ccr
      -- CP-element group 106: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Update/$entry
      -- 
    ccr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(106), ack => call_stmt_1955_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "ReceiveEngineDaemon_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_3116_elements(108);
      gj_ReceiveEngineDaemon_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	66 
    -- CP-element group 107: 	54 
    -- CP-element group 107: 	102 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Sample/cra
      -- CP-element group 107: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Sample/$exit
      -- 
    cra_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1955_call_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(107)); -- 
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	116 
    -- CP-element group 108: 	109 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	35 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/ring_reenable_memory_space_0
      -- CP-element group 108: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_Update/cca
      -- CP-element group 108: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1955_update_completed_
      -- 
    cca_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1955_call_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	100 
    -- CP-element group 109: 	104 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/barrier_stmt_1956_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Sample/req
      -- CP-element group 109: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_sample_start_
      -- 
    req_3551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(109), ack => WPIPE_RX_ACTIVITY_LOGGER_1957_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 3);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "ReceiveEngineDaemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(100) & ReceiveEngineDaemon_CP_3116_elements(104) & ReceiveEngineDaemon_CP_3116_elements(108);
      gj_ReceiveEngineDaemon_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Sample/ack
      -- CP-element group 110: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Update/req
      -- 
    ack_3552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1957_inst_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(110)); -- 
    req_3556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(110), ack => WPIPE_RX_ACTIVITY_LOGGER_1957_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	116 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	39 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Update/ack
      -- CP-element group 111: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/WPIPE_RX_ACTIVITY_LOGGER_1957_update_completed_
      -- 
    ack_3557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_RX_ACTIVITY_LOGGER_1957_inst_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(111)); -- 
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	14 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	15 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(14), ack => ReceiveEngineDaemon_CP_3116_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	38 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	85 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1839_call_stmt_1923_delay
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(113) is a control-delay.
    cp_element_113_delay: control_delay_element  generic map(name => " 113_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(38), ack => ReceiveEngineDaemon_CP_3116_elements(113), clk => clk, reset =>reset);
    -- CP-element group 114:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	88 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	93 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1923_call_stmt_1939_delay
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(114) is a control-delay.
    cp_element_114_delay: control_delay_element  generic map(name => " 114_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(88), ack => ReceiveEngineDaemon_CP_3116_elements(114), clk => clk, reset =>reset);
    -- CP-element group 115:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	96 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	105 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/call_stmt_1939_call_stmt_1955_delay
      -- 
    -- Element group ReceiveEngineDaemon_CP_3116_elements(115) is a control-delay.
    cp_element_115_delay: control_delay_element  generic map(name => " 115_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_3116_elements(96), ack => ReceiveEngineDaemon_CP_3116_elements(115), clk => clk, reset =>reset);
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	111 
    -- CP-element group 116: 	108 
    -- CP-element group 116: 	17 
    -- CP-element group 116: 	20 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	11 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1812/do_while_stmt_1825/do_while_stmt_1825_loop_body/$exit
      -- 
    ReceiveEngineDaemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 3,1 => 3,2 => 3,3 => 3);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "ReceiveEngineDaemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_3116_elements(111) & ReceiveEngineDaemon_CP_3116_elements(108) & ReceiveEngineDaemon_CP_3116_elements(17) & ReceiveEngineDaemon_CP_3116_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	10 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_exit/ack
      -- CP-element group 117: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_exit/$exit
      -- 
    ack_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1825_branch_ack_0, ack => ReceiveEngineDaemon_CP_3116_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	10 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_taken/$exit
      -- CP-element group 118: 	 branch_block_stmt_1812/do_while_stmt_1825/loop_taken/ack
      -- 
    ack_3570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1825_branch_ack_1, ack => ReceiveEngineDaemon_CP_3116_elements(118)); -- 
    -- CP-element group 119:  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	8 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	4 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1812/do_while_stmt_1825/$exit
      -- 
    ReceiveEngineDaemon_CP_3116_elements(119) <= ReceiveEngineDaemon_CP_3116_elements(8);
    -- CP-element group 120:  merge  branch  transition  place  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	2 
    -- CP-element group 120: 	4 
    -- CP-element group 120: 	5 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	5 
    -- CP-element group 120: 	6 
    -- CP-element group 120:  members (49) 
      -- CP-element group 120: 	 branch_block_stmt_1812/merge_stmt_1813_PhiReqMerge
      -- CP-element group 120: 	 branch_block_stmt_1812/merge_stmt_1813__exit__
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814__entry__
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_dead_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Sample/req
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Update/req
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_S_CONTROL_REGISTER_1815/Update/ack
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/cr
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/cr
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_eval_test/branch_req
      -- CP-element group 120: 	 branch_block_stmt_1812/NOT_u1_u1_1818_place
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_if_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/if_stmt_1814_else_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/merge_stmt_1813_PhiAck/$entry
      -- CP-element group 120: 	 branch_block_stmt_1812/merge_stmt_1813_PhiAck/$exit
      -- CP-element group 120: 	 branch_block_stmt_1812/merge_stmt_1813_PhiAck/dummy
      -- 
    branch_req_3205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_3116_elements(120), ack => if_stmt_1814_branch_req_0); -- 
    ReceiveEngineDaemon_CP_3116_elements(120) <= OrReduce(ReceiveEngineDaemon_CP_3116_elements(2) & ReceiveEngineDaemon_CP_3116_elements(4) & ReceiveEngineDaemon_CP_3116_elements(5));
    ReceiveEngineDaemon_do_while_stmt_1825_terminator_3571: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_1825_terminator_3571", max_iterations_in_flight =>3) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_3116_elements(11),loop_continue => ReceiveEngineDaemon_CP_3116_elements(118),loop_terminate => ReceiveEngineDaemon_CP_3116_elements(117),loop_back => ReceiveEngineDaemon_CP_3116_elements(9),loop_exit => ReceiveEngineDaemon_CP_3116_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1827_phi_seq_3273_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ReceiveEngineDaemon_CP_3116_elements(22);
      ReceiveEngineDaemon_CP_3116_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ReceiveEngineDaemon_CP_3116_elements(27);
      ReceiveEngineDaemon_CP_3116_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= ReceiveEngineDaemon_CP_3116_elements(29);
      ReceiveEngineDaemon_CP_3116_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= ReceiveEngineDaemon_CP_3116_elements(24);
      ReceiveEngineDaemon_CP_3116_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ReceiveEngineDaemon_CP_3116_elements(31);
      ReceiveEngineDaemon_CP_3116_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= ReceiveEngineDaemon_CP_3116_elements(33);
      ReceiveEngineDaemon_CP_3116_elements(25) <= phi_mux_reqs(1);
      phi_stmt_1827_phi_seq_3273 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_1827_phi_seq_3273") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ReceiveEngineDaemon_CP_3116_elements(16), 
          phi_sample_ack => ReceiveEngineDaemon_CP_3116_elements(20), 
          phi_update_req => ReceiveEngineDaemon_CP_3116_elements(19), 
          phi_update_ack => ReceiveEngineDaemon_CP_3116_elements(21), 
          phi_mux_ack => ReceiveEngineDaemon_CP_3116_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3234_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_3116_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_3116_elements(13);
        entry_tmerge_3234 : transition_merge -- 
          generic map(name => " entry_tmerge_3234")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_3116_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1800_1800_delayed_43_0_1897 : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_1817_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1964_wire : std_logic_vector(0 downto 0);
    signal MUX_1908_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_1781_1781_delayed_39_0_1876 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1788_1788_delayed_39_0_1886 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1818_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1880_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1919_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_S_CONTROL_REGISTER_1815_wire : std_logic_vector(31 downto 0);
    signal RPIPE_S_CONTROL_REGISTER_1962_wire : std_logic_vector(31 downto 0);
    signal R_FREEQUEUE_1835_wire_constant : std_logic_vector(1 downto 0);
    signal R_FREEQUEUE_1951_wire_constant : std_logic_vector(1 downto 0);
    signal R_READMEM_1845_wire_constant : std_logic_vector(0 downto 0);
    signal bad_packet_identifier_1868 : std_logic_vector(0 downto 0);
    signal cond_1928 : std_logic_vector(0 downto 0);
    signal control_dword_1852 : std_logic_vector(63 downto 0);
    signal free_flag_1891 : std_logic_vector(0 downto 0);
    signal ignore_resp1_1923 : std_logic_vector(31 downto 0);
    signal init_flag_1793_delayed_42_0_1900 : std_logic_vector(0 downto 0);
    signal init_flag_1827 : std_logic_vector(0 downto 0);
    signal konst_1810_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1816_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1836_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1871_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1920_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1926_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1942_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1952_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1958_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1963_wire_constant : std_logic_vector(31 downto 0);
    signal max_buffer_addr_offset_1856 : std_logic_vector(15 downto 0);
    signal ok_flag_1805_delayed_1_0_1913 : std_logic_vector(0 downto 0);
    signal ok_flag_1882 : std_logic_vector(0 downto 0);
    signal pkt_cnt_1910 : std_logic_vector(31 downto 0);
    signal push_status_1955 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_1772_delayed_38_0_1862 : std_logic_vector(63 downto 0);
    signal rx_buffer_pointer_1826_delayed_39_0_1935 : std_logic_vector(63 downto 0);
    signal rx_buffer_pointer_1838_delayed_39_0_1948 : std_logic_vector(63 downto 0);
    signal rx_buffer_pointer_1839 : std_logic_vector(63 downto 0);
    signal rx_tag_1824 : std_logic_vector(7 downto 0);
    signal status_1769_delayed_38_0_1859 : std_logic_vector(0 downto 0);
    signal status_1839 : std_logic_vector(0 downto 0);
    signal type_cast_1830_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1832_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1848_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1850_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1895_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1904_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1916_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1919_wire_constant <= "1111";
    R_FREEQUEUE_1835_wire_constant <= "00";
    R_FREEQUEUE_1951_wire_constant <= "00";
    R_READMEM_1845_wire_constant <= "1";
    konst_1810_wire_constant <= "00000000";
    konst_1816_wire_constant <= "00000000000000000000000000000000";
    konst_1836_wire_constant <= "00000000";
    konst_1841_wire_constant <= "00000001";
    konst_1871_wire_constant <= "00000010";
    konst_1920_wire_constant <= "00000011";
    konst_1926_wire_constant <= "1";
    konst_1942_wire_constant <= "00000011";
    konst_1952_wire_constant <= "00000000";
    konst_1958_wire_constant <= "00000100";
    konst_1963_wire_constant <= "00000000000000000000000000000000";
    rx_tag_1824 <= "00000001";
    type_cast_1830_wire_constant <= "0";
    type_cast_1832_wire_constant <= "1";
    type_cast_1848_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1850_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1895_wire_constant <= "00000000000000000000000000000001";
    type_cast_1904_wire_constant <= "00000000000000000000000000000001";
    type_cast_1916_wire_constant <= "0";
    phi_stmt_1827: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1830_wire_constant & type_cast_1832_wire_constant;
      req <= phi_stmt_1827_req_0 & phi_stmt_1827_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1827",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1827_ack_0,
          idata => idata,
          odata => init_flag_1827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1827
    -- flow-through select operator MUX_1908_inst
    MUX_1908_wire <= ADD_u32_u32_1800_1800_delayed_43_0_1897 when (ok_flag_1882(0) /=  '0') else pkt_cnt_1910;
    MUX_1909_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1909_inst_req_0;
      MUX_1909_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1909_inst_req_1;
      MUX_1909_inst_ack_1<= update_ack(0);
      MUX_1909_inst: SelectSplitProtocol generic map(name => "MUX_1909_inst", data_width => 32, buffering => 2, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_1904_wire_constant, y => MUX_1908_wire, sel => init_flag_1793_delayed_42_0_1900, z => pkt_cnt_1910, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_1855_inst
    max_buffer_addr_offset_1856 <= control_dword_1852(63 downto 48);
    W_init_flag_1793_delayed_42_0_1898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_init_flag_1793_delayed_42_0_1898_inst_req_0;
      W_init_flag_1793_delayed_42_0_1898_inst_ack_0<= wack(0);
      rreq(0) <= W_init_flag_1793_delayed_42_0_1898_inst_req_1;
      W_init_flag_1793_delayed_42_0_1898_inst_ack_1<= rack(0);
      W_init_flag_1793_delayed_42_0_1898_inst : InterlockBuffer generic map ( -- 
        name => "W_init_flag_1793_delayed_42_0_1898_inst",
        buffer_size => 42,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => init_flag_1827,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => init_flag_1793_delayed_42_0_1900,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ok_flag_1805_delayed_1_0_1911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ok_flag_1805_delayed_1_0_1911_inst_req_0;
      W_ok_flag_1805_delayed_1_0_1911_inst_ack_0<= wack(0);
      rreq(0) <= W_ok_flag_1805_delayed_1_0_1911_inst_req_1;
      W_ok_flag_1805_delayed_1_0_1911_inst_ack_1<= rack(0);
      W_ok_flag_1805_delayed_1_0_1911_inst : InterlockBuffer generic map ( -- 
        name => "W_ok_flag_1805_delayed_1_0_1911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ok_flag_1882,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ok_flag_1805_delayed_1_0_1913,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_req_0;
      W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_req_1;
      W_rx_buffer_pointer_1772_delayed_38_0_1860_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1772_delayed_38_0_1860_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1772_delayed_38_0_1860_inst",
        buffer_size => 38,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_1839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1772_delayed_38_0_1862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_req_0;
      W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_req_1;
      W_rx_buffer_pointer_1826_delayed_39_0_1933_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1826_delayed_39_0_1933_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1826_delayed_39_0_1933_inst",
        buffer_size => 39,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_1839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1826_delayed_39_0_1935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_req_0;
      W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_req_1;
      W_rx_buffer_pointer_1838_delayed_39_0_1946_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1838_delayed_39_0_1946_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1838_delayed_39_0_1946_inst",
        buffer_size => 39,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_1839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1838_delayed_39_0_1948,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_status_1769_delayed_38_0_1857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_1769_delayed_38_0_1857_inst_req_0;
      W_status_1769_delayed_38_0_1857_inst_ack_0<= wack(0);
      rreq(0) <= W_status_1769_delayed_38_0_1857_inst_req_1;
      W_status_1769_delayed_38_0_1857_inst_ack_1<= rack(0);
      W_status_1769_delayed_38_0_1857_inst : InterlockBuffer generic map ( -- 
        name => "W_status_1769_delayed_38_0_1857_inst",
        buffer_size => 38,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => status_1839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_1769_delayed_38_0_1859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1825_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1964_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1825_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1825_branch_req_0,
          ack0 => do_while_stmt_1825_branch_ack_0,
          ack1 => do_while_stmt_1825_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1814_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1818_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1814_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1814_branch_req_0,
          ack0 => if_stmt_1814_branch_ack_0,
          ack1 => if_stmt_1814_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_1896_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 43);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pkt_cnt_1910;
      ADD_u32_u32_1800_1800_delayed_43_0_1897 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_1896_inst_req_0;
      ADD_u32_u32_1896_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_1896_inst_req_1;
      ADD_u32_u32_1896_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 43,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- flow through binary operator AND_u1_u1_1881_inst
    ok_flag_1882 <= (NOT_u1_u1_1781_1781_delayed_39_0_1876 and NOT_u1_u1_1880_wire);
    -- flow through binary operator AND_u1_u1_1890_inst
    free_flag_1891 <= (NOT_u1_u1_1788_1788_delayed_39_0_1886 and bad_packet_identifier_1868);
    -- flow through binary operator BITSEL_u32_u1_1817_inst
    process(RPIPE_S_CONTROL_REGISTER_1815_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_S_CONTROL_REGISTER_1815_wire, konst_1816_wire_constant, tmp_var);
      BITSEL_u32_u1_1817_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_1964_inst
    process(RPIPE_S_CONTROL_REGISTER_1962_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_S_CONTROL_REGISTER_1962_wire, konst_1963_wire_constant, tmp_var);
      BITSEL_u32_u1_1964_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_1927_inst
    process(ok_flag_1882) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ok_flag_1882, konst_1926_wire_constant, tmp_var);
      cond_1928 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1818_inst
    process(BITSEL_u32_u1_1817_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1817_wire, tmp_var);
      NOT_u1_u1_1818_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (7) : NOT_u1_u1_1875_inst 
    ApIntNot_group_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 39);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1839;
      NOT_u1_u1_1781_1781_delayed_39_0_1876 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1875_inst_req_0;
      NOT_u1_u1_1875_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1875_inst_req_1;
      NOT_u1_u1_1875_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_7_gI: SplitGuardInterface generic map(name => "ApIntNot_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 39,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- unary operator NOT_u1_u1_1880_inst
    process(bad_packet_identifier_1868) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_1868, tmp_var);
      NOT_u1_u1_1880_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (9) : NOT_u1_u1_1885_inst 
    ApIntNot_group_9: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 39);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1839;
      NOT_u1_u1_1788_1788_delayed_39_0_1886 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1885_inst_req_0;
      NOT_u1_u1_1885_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1885_inst_req_1;
      NOT_u1_u1_1885_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_9_gI: SplitGuardInterface generic map(name => "ApIntNot_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 39,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- read from input-signal S_CONTROL_REGISTER
    RPIPE_S_CONTROL_REGISTER_1815_wire <= S_CONTROL_REGISTER;
    RPIPE_S_CONTROL_REGISTER_1962_wire <= S_CONTROL_REGISTER;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1809_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1810_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_RX_ACTIVITY_LOGGER_1840_inst WPIPE_RX_ACTIVITY_LOGGER_1870_inst WPIPE_RX_ACTIVITY_LOGGER_1941_inst WPIPE_RX_ACTIVITY_LOGGER_1957_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_RX_ACTIVITY_LOGGER_1840_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_RX_ACTIVITY_LOGGER_1870_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_RX_ACTIVITY_LOGGER_1941_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_RX_ACTIVITY_LOGGER_1957_inst_req_0;
      WPIPE_RX_ACTIVITY_LOGGER_1840_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_RX_ACTIVITY_LOGGER_1870_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_RX_ACTIVITY_LOGGER_1941_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_RX_ACTIVITY_LOGGER_1957_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_RX_ACTIVITY_LOGGER_1840_inst_req_1;
      update_req_unguarded(2) <= WPIPE_RX_ACTIVITY_LOGGER_1870_inst_req_1;
      update_req_unguarded(1) <= WPIPE_RX_ACTIVITY_LOGGER_1941_inst_req_1;
      update_req_unguarded(0) <= WPIPE_RX_ACTIVITY_LOGGER_1957_inst_req_1;
      WPIPE_RX_ACTIVITY_LOGGER_1840_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_RX_ACTIVITY_LOGGER_1870_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_RX_ACTIVITY_LOGGER_1941_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_RX_ACTIVITY_LOGGER_1957_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      data_in <= konst_1841_wire_constant & konst_1871_wire_constant & konst_1942_wire_constant & konst_1958_wire_constant;
      RX_ACTIVITY_LOGGER_write_1_gI: SplitGuardInterface generic map(name => "RX_ACTIVITY_LOGGER_write_1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      RX_ACTIVITY_LOGGER_write_1: OutputPortRevised -- 
        generic map ( name => "RX_ACTIVITY_LOGGER", data_width => 8, num_reqs => 4, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => RX_ACTIVITY_LOGGER_pipe_write_req(0),
          oack => RX_ACTIVITY_LOGGER_pipe_write_ack(0),
          odata => RX_ACTIVITY_LOGGER_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1839_call 
    popFromQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1839_call_req_0;
      call_stmt_1839_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1839_call_req_1;
      call_stmt_1839_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_0_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_tag_1824 & R_FREEQUEUE_1835_wire_constant & konst_1836_wire_constant;
      rx_buffer_pointer_1839 <= data_out(64 downto 1);
      status_1839 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 18,
        owidth => 18,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(17 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 65,
          owidth => 65,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(64 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1852_call 
    accessMemoryDword_call_group_1: Block -- 
      signal data_in: std_logic_vector(200 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 38);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1852_call_req_0;
      call_stmt_1852_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1852_call_req_1;
      call_stmt_1852_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDword_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_tag_1824 & R_READMEM_1845_wire_constant & rx_buffer_pointer_1839 & type_cast_1848_wire_constant & type_cast_1850_wire_constant;
      control_dword_1852 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 201,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(0),
          ackR => accessMemoryDword_call_acks(0),
          dataR => accessMemoryDword_call_data(200 downto 0),
          tagR => accessMemoryDword_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(0), -- cross-over
          ackL => accessMemoryDword_return_reqs(0), -- cross-over
          dataL => accessMemoryDword_return_data(63 downto 0),
          tagL => accessMemoryDword_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1868_call 
    loadBuffer_call_group_2: Block -- 
      signal data_in: std_logic_vector(87 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1868_call_req_0;
      call_stmt_1868_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1868_call_req_1;
      call_stmt_1868_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_1769_delayed_38_0_1859(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_2_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_tag_1824 & max_buffer_addr_offset_1856 & rx_buffer_pointer_1772_delayed_38_0_1862;
      bad_packet_identifier_1868 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 88,
        owidth => 88,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(87 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1923_call 
    accessRegister_call_group_3: Block -- 
      signal data_in: std_logic_vector(44 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1923_call_req_0;
      call_stmt_1923_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1923_call_req_1;
      call_stmt_1923_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1805_delayed_1_0_1913(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessRegister_call_group_3_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1916_wire_constant & NOT_u4_u4_1919_wire_constant & konst_1920_wire_constant & pkt_cnt_1910;
      ignore_resp1_1923 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 45,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1939_call 
    populateRxQueue_call_group_4: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1939_call_req_0;
      call_stmt_1939_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1939_call_req_1;
      call_stmt_1939_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1882(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_4_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_tag_1824 & rx_buffer_pointer_1826_delayed_39_0_1935;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(71 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1955_call 
    pushIntoQueue_call_group_5: Block -- 
      signal data_in: std_logic_vector(81 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1955_call_req_0;
      call_stmt_1955_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1955_call_req_1;
      call_stmt_1955_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_1891(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_5_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_tag_1824 & R_FREEQUEUE_1951_wire_constant & konst_1952_wire_constant & rx_buffer_pointer_1838_delayed_39_0_1948;
      push_status_1955 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 82,
        owidth => 82,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(81 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryBase is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    request : in  std_logic_vector(109 downto 0);
    response : out  std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_DEBUG_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_DEBUG_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_DEBUG_SIGNAL_pipe_write_data : out  std_logic_vector(255 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryBase;
architecture accessMemoryBase_arch of accessMemoryBase is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 118)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 65)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal request_buffer :  std_logic_vector(109 downto 0);
  signal request_update_enable: Boolean;
  -- output port buffer signals
  signal response_buffer :  std_logic_vector(64 downto 0);
  signal response_update_enable: Boolean;
  signal accessMemoryBase_CP_226_start: Boolean;
  signal accessMemoryBase_CP_226_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_DEBUG_SIGNAL_306_inst_req_0 : boolean;
  signal WPIPE_NIC_DEBUG_SIGNAL_306_inst_ack_0 : boolean;
  signal WPIPE_NIC_DEBUG_SIGNAL_306_inst_req_1 : boolean;
  signal WPIPE_NIC_DEBUG_SIGNAL_306_inst_ack_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_ack_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryBase_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 118) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(117 downto 8) <= request;
  request_buffer <= in_buffer_data_out(117 downto 8);
  in_buffer_data_in(tag_length + 117 downto 118) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 117 downto 118);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 1,3 => 7);
    constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 7);
    constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 4); -- 
  begin -- 
    preds <= tag_update_enable & request_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryBase_CP_226_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryBase_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 65) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(64 downto 0) <= response_buffer;
  response <= out_buffer_data_out(64 downto 0);
  out_buffer_data_in(tag_length + 64 downto 65) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 64 downto 65);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryBase_CP_226_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  response_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 27) := "response_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_response_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => response_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryBase_CP_226_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryBase_CP_226_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryBase_CP_226: Block -- control-path 
    signal accessMemoryBase_CP_226_elements: BooleanArray(19 downto 0);
    -- 
  begin -- 
    accessMemoryBase_CP_226_elements(0) <= accessMemoryBase_CP_226_start;
    accessMemoryBase_CP_226_symbol <= accessMemoryBase_CP_226_elements(19);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	12 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_292_to_assign_stmt_308/$entry
      -- 
    accessMemoryBase_CP_226_elements(1) <= accessMemoryBase_CP_226_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	13 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_292_to_assign_stmt_308/tag_update_enable
      -- CP-element group 2: 	 assign_stmt_292_to_assign_stmt_308/tag_update_enable_out
      -- 
    accessMemoryBase_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryBase_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryBase_CP_226_elements(13);
      gj_accessMemoryBase_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	6 
    -- CP-element group 3: 	13 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_292_to_assign_stmt_308/request_update_enable
      -- CP-element group 3: 	 assign_stmt_292_to_assign_stmt_308/request_update_enable_out
      -- 
    accessMemoryBase_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "accessMemoryBase_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryBase_CP_226_elements(6) & accessMemoryBase_CP_226_elements(13);
      gj_accessMemoryBase_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	9 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_292_to_assign_stmt_308/response_update_enable
      -- CP-element group 4: 	 assign_stmt_292_to_assign_stmt_308/response_update_enable_in
      -- 
    accessMemoryBase_CP_226_elements(4) <= accessMemoryBase_CP_226_elements(18);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_sample_start_
      -- CP-element group 5: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Sample/req
      -- 
    req_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryBase_CP_226_elements(5), ack => WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_req_0); -- 
    accessMemoryBase_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "accessMemoryBase_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryBase_CP_226_elements(1) & accessMemoryBase_CP_226_elements(7);
      gj_accessMemoryBase_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	3 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_sample_completed_
      -- CP-element group 6: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_update_start_
      -- CP-element group 6: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Sample/ack
      -- CP-element group 6: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Update/$entry
      -- CP-element group 6: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Update/req
      -- 
    ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_ack_0, ack => accessMemoryBase_CP_226_elements(6)); -- 
    req_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryBase_CP_226_elements(6), ack => WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	15 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_update_completed_
      -- CP-element group 7: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Update/$exit
      -- CP-element group 7: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_TO_MEMORY_REQUEST_290_Update/ack
      -- 
    ack_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_ack_1, ack => accessMemoryBase_CP_226_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	11 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_sample_start_
      -- CP-element group 8: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Sample/rr
      -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryBase_CP_226_elements(8), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_req_0); -- 
    accessMemoryBase_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "accessMemoryBase_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryBase_CP_226_elements(1) & accessMemoryBase_CP_226_elements(11);
      gj_accessMemoryBase_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	4 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_update_start_
      -- CP-element group 9: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Update/$entry
      -- CP-element group 9: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Update/cr
      -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryBase_CP_226_elements(9), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_req_1); -- 
    accessMemoryBase_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "accessMemoryBase_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMemoryBase_CP_226_elements(10) & accessMemoryBase_CP_226_elements(4) & accessMemoryBase_CP_226_elements(13);
      gj_accessMemoryBase_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	9 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_sample_completed_
      -- CP-element group 10: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Sample/$exit
      -- CP-element group 10: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_ack_0, ack => accessMemoryBase_CP_226_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	8 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_update_completed_
      -- CP-element group 11: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Update/$exit
      -- CP-element group 11: 	 assign_stmt_292_to_assign_stmt_308/RPIPE_MEMORY_TO_NIC_RESPONSE_294_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_ack_1, ack => accessMemoryBase_CP_226_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: 	1 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_sample_start_
      -- CP-element group 12: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Sample/$entry
      -- CP-element group 12: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Sample/req
      -- 
    req_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryBase_CP_226_elements(12), ack => WPIPE_NIC_DEBUG_SIGNAL_306_inst_req_0); -- 
    accessMemoryBase_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "accessMemoryBase_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMemoryBase_CP_226_elements(11) & accessMemoryBase_CP_226_elements(1) & accessMemoryBase_CP_226_elements(14);
      gj_accessMemoryBase_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: 	2 
    -- CP-element group 13: 	3 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_sample_completed_
      -- CP-element group 13: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_update_start_
      -- CP-element group 13: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Sample/ack
      -- CP-element group 13: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Update/$entry
      -- CP-element group 13: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Update/req
      -- 
    ack_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_DEBUG_SIGNAL_306_inst_ack_0, ack => accessMemoryBase_CP_226_elements(13)); -- 
    req_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryBase_CP_226_elements(13), ack => WPIPE_NIC_DEBUG_SIGNAL_306_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_update_completed_
      -- CP-element group 14: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Update/$exit
      -- CP-element group 14: 	 assign_stmt_292_to_assign_stmt_308/WPIPE_NIC_DEBUG_SIGNAL_306_Update/ack
      -- 
    ack_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_DEBUG_SIGNAL_306_inst_ack_1, ack => accessMemoryBase_CP_226_elements(14)); -- 
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	7 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	19 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_292_to_assign_stmt_308/$exit
      -- 
    accessMemoryBase_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "accessMemoryBase_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryBase_CP_226_elements(7) & accessMemoryBase_CP_226_elements(14);
      gj_accessMemoryBase_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryBase_CP_226_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 tag_update_enable
      -- 
    accessMemoryBase_CP_226_elements(16) <= accessMemoryBase_CP_226_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 request_update_enable
      -- 
    accessMemoryBase_CP_226_elements(17) <= accessMemoryBase_CP_226_elements(3);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 response_update_enable
      -- 
    -- CP-element group 19:  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 $exit
      -- 
    accessMemoryBase_CP_226_elements(19) <= accessMemoryBase_CP_226_elements(15);
    --  hookup: inputs to control-path 
    accessMemoryBase_CP_226_elements(18) <= response_update_enable;
    -- hookup: output from control-path 
    tag_update_enable <= accessMemoryBase_CP_226_elements(16);
    request_update_enable <= accessMemoryBase_CP_226_elements(17);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u110_u175_303_wire : std_logic_vector(174 downto 0);
    signal CONCAT_u73_u81_300_wire : std_logic_vector(80 downto 0);
    signal debug_sig_305 : std_logic_vector(255 downto 0);
    signal type_cast_298_wire_constant : std_logic_vector(72 downto 0);
    -- 
  begin -- 
    type_cast_298_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000";
    -- flow through binary operator CONCAT_u110_u175_303_inst
    process(request_buffer, response_buffer) -- 
      variable tmp_var : std_logic_vector(174 downto 0); -- 
    begin -- 
      ApConcat_proc(request_buffer, response_buffer, tmp_var);
      CONCAT_u110_u175_303_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u73_u81_300_inst
    process(type_cast_298_wire_constant, tag_buffer) -- 
      variable tmp_var : std_logic_vector(80 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_298_wire_constant, tag_buffer, tmp_var);
      CONCAT_u73_u81_300_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u81_u256_304_inst
    process(CONCAT_u73_u81_300_wire, CONCAT_u110_u175_303_wire) -- 
      variable tmp_var : std_logic_vector(255 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u73_u81_300_wire, CONCAT_u110_u175_303_wire, tmp_var);
      debug_sig_305 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_294_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_buffer <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_DEBUG_SIGNAL_306_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_DEBUG_SIGNAL_306_inst_req_0;
      WPIPE_NIC_DEBUG_SIGNAL_306_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_DEBUG_SIGNAL_306_inst_req_1;
      WPIPE_NIC_DEBUG_SIGNAL_306_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= debug_sig_305;
      NIC_DEBUG_SIGNAL_write_0_gI: SplitGuardInterface generic map(name => "NIC_DEBUG_SIGNAL_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_DEBUG_SIGNAL_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_DEBUG_SIGNAL", data_width => 256, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_DEBUG_SIGNAL_pipe_write_req(0),
          oack => NIC_DEBUG_SIGNAL_pipe_write_ack(0),
          odata => NIC_DEBUG_SIGNAL_pipe_write_data(255 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_NIC_TO_MEMORY_REQUEST_290_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_290_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_buffer;
      NIC_TO_MEMORY_REQUEST_write_1_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_1: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end accessMemoryBase_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryByte is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    byte_addr_base : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wbyte : in  std_logic_vector(7 downto 0);
    rbyte : out  std_logic_vector(7 downto 0);
    doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_call_data : out  std_logic_vector(202 downto 0);
    doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
    doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_return_data : in   std_logic_vector(63 downto 0);
    doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryByte;
architecture accessMemoryByte_arch of accessMemoryByte is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 145)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal byte_addr_base_buffer :  std_logic_vector(63 downto 0);
  signal byte_addr_base_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wbyte_buffer :  std_logic_vector(7 downto 0);
  signal wbyte_update_enable: Boolean;
  -- output port buffer signals
  signal rbyte_buffer :  std_logic_vector(7 downto 0);
  signal rbyte_update_enable: Boolean;
  signal accessMemoryByte_CP_1611_start: Boolean;
  signal accessMemoryByte_CP_1611_symbol: Boolean;
  -- volatile/operator module components. 
  component doMemAccess is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      opcode : in  std_logic_vector(2 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      memory_access_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_data : out  std_logic_vector(169 downto 0);
      accessMemoryWordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWordBase_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_data : out  std_logic_vector(145 downto 0);
      accessMemoryByteBase_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryByteBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByteBase_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemoryDwordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_data : out  std_logic_vector(201 downto 0);
      accessMemoryDwordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDwordBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1182_call_req_1 : boolean;
  signal call_stmt_1182_call_req_0 : boolean;
  signal call_stmt_1182_call_ack_1 : boolean;
  signal call_stmt_1182_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryByte_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 145) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= byte_addr_base;
  byte_addr_base_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(136 downto 73) <= offset;
  offset_buffer <= in_buffer_data_out(136 downto 73);
  in_buffer_data_in(144 downto 137) <= wbyte;
  wbyte_buffer <= in_buffer_data_out(144 downto 137);
  in_buffer_data_in(tag_length + 144 downto 145) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 144 downto 145);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 1,6 => 7);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 7);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= tag_update_enable & rwbar_update_enable & byte_addr_base_update_enable & offset_update_enable & wbyte_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryByte_CP_1611_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryByte_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= rbyte_buffer;
  rbyte <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryByte_CP_1611_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rbyte_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rbyte_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rbyte_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rbyte_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryByte_CP_1611_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryByte_CP_1611_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryByte_CP_1611: Block -- control-path 
    signal accessMemoryByte_CP_1611_elements: BooleanArray(18 downto 0);
    -- 
  begin -- 
    accessMemoryByte_CP_1611_elements(0) <= accessMemoryByte_CP_1611_start;
    accessMemoryByte_CP_1611_symbol <= accessMemoryByte_CP_1611_elements(18);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1182_to_assign_stmt_1186/$entry
      -- 
    accessMemoryByte_CP_1611_elements(1) <= accessMemoryByte_CP_1611_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1182_to_assign_stmt_1186/tag_update_enable_out
      -- CP-element group 2: 	 call_stmt_1182_to_assign_stmt_1186/tag_update_enable
      -- 
    accessMemoryByte_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByte_CP_1611_elements(10);
      gj_accessMemoryByte_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	10 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1182_to_assign_stmt_1186/rwbar_update_enable
      -- CP-element group 3: 	 call_stmt_1182_to_assign_stmt_1186/rwbar_update_enable_out
      -- 
    accessMemoryByte_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByte_CP_1611_elements(10);
      gj_accessMemoryByte_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	10 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	14 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_1182_to_assign_stmt_1186/byte_addr_base_update_enable
      -- CP-element group 4: 	 call_stmt_1182_to_assign_stmt_1186/byte_addr_base_update_enable_out
      -- 
    accessMemoryByte_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByte_CP_1611_elements(10);
      gj_accessMemoryByte_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	15 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_1182_to_assign_stmt_1186/offset_update_enable
      -- CP-element group 5: 	 call_stmt_1182_to_assign_stmt_1186/offset_update_enable_out
      -- 
    accessMemoryByte_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByte_CP_1611_elements(10);
      gj_accessMemoryByte_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	10 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	16 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 call_stmt_1182_to_assign_stmt_1186/wbyte_update_enable_out
      -- CP-element group 6: 	 call_stmt_1182_to_assign_stmt_1186/wbyte_update_enable
      -- 
    accessMemoryByte_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByte_CP_1611_elements(10);
      gj_accessMemoryByte_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	17 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 call_stmt_1182_to_assign_stmt_1186/rbyte_update_enable
      -- CP-element group 7: 	 call_stmt_1182_to_assign_stmt_1186/rbyte_update_enable_in
      -- 
    accessMemoryByte_CP_1611_elements(7) <= accessMemoryByte_CP_1611_elements(17);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_sample_start_
      -- CP-element group 8: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Sample/crr
      -- 
    crr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByte_CP_1611_elements(8), ack => call_stmt_1182_call_req_0); -- 
    accessMemoryByte_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByte_CP_1611_elements(1) & accessMemoryByte_CP_1611_elements(10);
      gj_accessMemoryByte_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Update/ccr
      -- CP-element group 9: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Update/$entry
      -- CP-element group 9: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_update_start_
      -- 
    ccr_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByte_CP_1611_elements(9), ack => call_stmt_1182_call_req_1); -- 
    accessMemoryByte_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "accessMemoryByte_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByte_CP_1611_elements(7) & accessMemoryByte_CP_1611_elements(11);
      gj_accessMemoryByte_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByte_CP_1611_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: 	5 
    -- CP-element group 10: 	6 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_sample_completed_
      -- CP-element group 10: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Sample/$exit
      -- CP-element group 10: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Sample/cra
      -- 
    cra_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1182_call_ack_0, ack => accessMemoryByte_CP_1611_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	18 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 call_stmt_1182_to_assign_stmt_1186/$exit
      -- CP-element group 11: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Update/cca
      -- CP-element group 11: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_Update/$exit
      -- CP-element group 11: 	 call_stmt_1182_to_assign_stmt_1186/call_stmt_1182_update_completed_
      -- 
    cca_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1182_call_ack_1, ack => accessMemoryByte_CP_1611_elements(11)); -- 
    -- CP-element group 12:  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 tag_update_enable
      -- 
    accessMemoryByte_CP_1611_elements(12) <= accessMemoryByte_CP_1611_elements(2);
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 rwbar_update_enable
      -- 
    accessMemoryByte_CP_1611_elements(13) <= accessMemoryByte_CP_1611_elements(3);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	4 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 byte_addr_base_update_enable
      -- 
    accessMemoryByte_CP_1611_elements(14) <= accessMemoryByte_CP_1611_elements(4);
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	5 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 offset_update_enable
      -- 
    accessMemoryByte_CP_1611_elements(15) <= accessMemoryByte_CP_1611_elements(5);
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	6 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 wbyte_update_enable
      -- 
    accessMemoryByte_CP_1611_elements(16) <= accessMemoryByte_CP_1611_elements(6);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	7 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rbyte_update_enable
      -- 
    -- CP-element group 18:  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 $exit
      -- 
    accessMemoryByte_CP_1611_elements(18) <= accessMemoryByte_CP_1611_elements(11);
    --  hookup: inputs to control-path 
    accessMemoryByte_CP_1611_elements(17) <= rbyte_update_enable;
    -- hookup: output from control-path 
    wbyte_update_enable <= accessMemoryByte_CP_1611_elements(16);
    offset_update_enable <= accessMemoryByte_CP_1611_elements(15);
    byte_addr_base_update_enable <= accessMemoryByte_CP_1611_elements(14);
    rwbar_update_enable <= accessMemoryByte_CP_1611_elements(13);
    tag_update_enable <= accessMemoryByte_CP_1611_elements(12);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u56_u64_1180_wire : std_logic_vector(63 downto 0);
    signal MUX_1174_wire : std_logic_vector(2 downto 0);
    signal R_LDB_1172_wire_constant : std_logic_vector(2 downto 0);
    signal R_STB_1173_wire_constant : std_logic_vector(2 downto 0);
    signal rdword_1182 : std_logic_vector(63 downto 0);
    signal type_cast_1178_wire_constant : std_logic_vector(55 downto 0);
    -- 
  begin -- 
    R_LDB_1172_wire_constant <= "110";
    R_STB_1173_wire_constant <= "011";
    type_cast_1178_wire_constant <= "00000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_1174_inst
    MUX_1174_wire <= R_LDB_1172_wire_constant when (rwbar_buffer(0) /=  '0') else R_STB_1173_wire_constant;
    -- flow-through slice operator slice_1185_inst
    rbyte_buffer <= rdword_1182(7 downto 0);
    -- flow through binary operator CONCAT_u56_u64_1180_inst
    process(type_cast_1178_wire_constant, wbyte_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1178_wire_constant, wbyte_buffer, tmp_var);
      CONCAT_u56_u64_1180_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1182_call 
    doMemAccess_call_group_0: Block -- 
      signal data_in: std_logic_vector(202 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 36);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1182_call_req_0;
      call_stmt_1182_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1182_call_req_1;
      call_stmt_1182_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      doMemAccess_call_group_0_gI: SplitGuardInterface generic map(name => "doMemAccess_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & MUX_1174_wire & byte_addr_base_buffer & offset_buffer & CONCAT_u56_u64_1180_wire;
      rdword_1182 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 203,
        owidth => 203,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => doMemAccess_call_reqs(0),
          ackR => doMemAccess_call_acks(0),
          dataR => doMemAccess_call_data(202 downto 0),
          tagR => doMemAccess_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => doMemAccess_return_acks(0), -- cross-over
          ackL => doMemAccess_return_reqs(0), -- cross-over
          dataL => doMemAccess_return_data(63 downto 0),
          tagL => doMemAccess_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemoryByte_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryByteBase is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    byte_addr_base : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wbyte : in  std_logic_vector(7 downto 0);
    rbyte : out  std_logic_vector(7 downto 0);
    calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
    calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
    calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
    calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
    calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
    calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
    calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
    calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
    accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
    accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryByteBase;
architecture accessMemoryByteBase_arch of accessMemoryByteBase is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 146)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal byte_addr_base_buffer :  std_logic_vector(63 downto 0);
  signal byte_addr_base_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wbyte_buffer :  std_logic_vector(7 downto 0);
  signal wbyte_update_enable: Boolean;
  -- output port buffer signals
  signal rbyte_buffer :  std_logic_vector(7 downto 0);
  signal rbyte_update_enable: Boolean;
  signal accessMemoryByteBase_CP_283_start: Boolean;
  signal accessMemoryByteBase_CP_283_symbol: Boolean;
  -- volatile/operator module components. 
  component calculateAddress36 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      addr : out  std_logic_vector(35 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      request : in  std_logic_vector(109 downto 0);
      response : out  std_logic_vector(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_data : out  std_logic_vector(255 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal EQ_u3_u1_438_inst_ack_0 : boolean;
  signal EQ_u3_u1_438_inst_req_0 : boolean;
  signal OR_u8_u8_489_inst_req_1 : boolean;
  signal EQ_u3_u1_448_inst_ack_0 : boolean;
  signal OR_u8_u8_489_inst_ack_0 : boolean;
  signal EQ_u3_u1_448_inst_req_0 : boolean;
  signal OR_u8_u8_489_inst_req_0 : boolean;
  signal EQ_u3_u1_448_inst_ack_1 : boolean;
  signal EQ_u3_u1_448_inst_req_1 : boolean;
  signal EQ_u3_u1_433_inst_ack_1 : boolean;
  signal EQ_u3_u1_428_inst_ack_0 : boolean;
  signal EQ_u3_u1_428_inst_req_0 : boolean;
  signal EQ_u3_u1_428_inst_ack_1 : boolean;
  signal EQ_u3_u1_438_inst_ack_1 : boolean;
  signal EQ_u3_u1_438_inst_req_1 : boolean;
  signal EQ_u3_u1_433_inst_ack_0 : boolean;
  signal EQ_u3_u1_433_inst_req_1 : boolean;
  signal EQ_u3_u1_428_inst_req_1 : boolean;
  signal EQ_u3_u1_433_inst_req_0 : boolean;
  signal OR_u8_u8_489_inst_ack_1 : boolean;
  signal EQ_u3_u1_443_inst_ack_1 : boolean;
  signal EQ_u3_u1_443_inst_req_1 : boolean;
  signal EQ_u3_u1_443_inst_ack_0 : boolean;
  signal EQ_u3_u1_443_inst_req_0 : boolean;
  signal call_calculateAddress36_expr_321_inst_req_0 : boolean;
  signal call_calculateAddress36_expr_321_inst_ack_0 : boolean;
  signal call_calculateAddress36_expr_321_inst_req_1 : boolean;
  signal call_calculateAddress36_expr_321_inst_ack_1 : boolean;
  signal CONCAT_u8_u64_346_inst_req_0 : boolean;
  signal CONCAT_u8_u64_346_inst_ack_0 : boolean;
  signal CONCAT_u8_u64_346_inst_req_1 : boolean;
  signal CONCAT_u8_u64_346_inst_ack_1 : boolean;
  signal CONCAT_u1_u2_360_inst_req_0 : boolean;
  signal CONCAT_u1_u2_360_inst_ack_0 : boolean;
  signal CONCAT_u1_u2_360_inst_req_1 : boolean;
  signal CONCAT_u1_u2_360_inst_ack_1 : boolean;
  signal W_tag_365_delayed_3_0_371_inst_req_0 : boolean;
  signal W_tag_365_delayed_3_0_371_inst_ack_0 : boolean;
  signal W_tag_365_delayed_3_0_371_inst_req_1 : boolean;
  signal W_tag_365_delayed_3_0_371_inst_ack_1 : boolean;
  signal call_stmt_377_call_req_0 : boolean;
  signal call_stmt_377_call_ack_0 : boolean;
  signal call_stmt_377_call_req_1 : boolean;
  signal call_stmt_377_call_ack_1 : boolean;
  signal EQ_u3_u1_413_inst_req_0 : boolean;
  signal EQ_u3_u1_413_inst_ack_0 : boolean;
  signal EQ_u3_u1_413_inst_req_1 : boolean;
  signal EQ_u3_u1_413_inst_ack_1 : boolean;
  signal EQ_u3_u1_418_inst_req_0 : boolean;
  signal EQ_u3_u1_418_inst_ack_0 : boolean;
  signal EQ_u3_u1_418_inst_req_1 : boolean;
  signal EQ_u3_u1_418_inst_ack_1 : boolean;
  signal EQ_u3_u1_423_inst_req_0 : boolean;
  signal EQ_u3_u1_423_inst_ack_0 : boolean;
  signal EQ_u3_u1_423_inst_req_1 : boolean;
  signal EQ_u3_u1_423_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryByteBase_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 146) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= lock;
  lock_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(9 downto 9) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(9 downto 9);
  in_buffer_data_in(73 downto 10) <= byte_addr_base;
  byte_addr_base_buffer <= in_buffer_data_out(73 downto 10);
  in_buffer_data_in(137 downto 74) <= offset;
  offset_buffer <= in_buffer_data_out(137 downto 74);
  in_buffer_data_in(145 downto 138) <= wbyte;
  wbyte_buffer <= in_buffer_data_out(145 downto 138);
  in_buffer_data_in(tag_length + 145 downto 146) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 145 downto 146);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 1,7 => 7);
    constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1,7 => 7);
    constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 8); -- 
  begin -- 
    preds <= tag_update_enable & lock_update_enable & rwbar_update_enable & byte_addr_base_update_enable & offset_update_enable & wbyte_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryByteBase_CP_283_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryByteBase_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= rbyte_buffer;
  rbyte <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryByteBase_CP_283_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rbyte_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rbyte_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rbyte_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rbyte_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryByteBase_CP_283_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryByteBase_CP_283_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryByteBase_CP_283: Block -- control-path 
    signal accessMemoryByteBase_CP_283_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    accessMemoryByteBase_CP_283_elements(0) <= accessMemoryByteBase_CP_283_start;
    accessMemoryByteBase_CP_283_symbol <= accessMemoryByteBase_CP_283_elements(72);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	21 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_322_to_assign_stmt_490/$entry
      -- 
    accessMemoryByteBase_CP_283_elements(1) <= accessMemoryByteBase_CP_283_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	23 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	65 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_322_to_assign_stmt_490/tag_update_enable
      -- CP-element group 2: 	 assign_stmt_322_to_assign_stmt_490/tag_update_enable_out
      -- 
    accessMemoryByteBase_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByteBase_CP_283_elements(23);
      gj_accessMemoryByteBase_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	19 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	66 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_490/lock_update_enable
      -- CP-element group 3: 	 assign_stmt_322_to_assign_stmt_490/lock_update_enable_out
      -- 
    accessMemoryByteBase_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByteBase_CP_283_elements(19);
      gj_accessMemoryByteBase_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	19 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	67 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_322_to_assign_stmt_490/rwbar_update_enable
      -- CP-element group 4: 	 assign_stmt_322_to_assign_stmt_490/rwbar_update_enable_out
      -- 
    accessMemoryByteBase_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByteBase_CP_283_elements(19);
      gj_accessMemoryByteBase_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	68 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_322_to_assign_stmt_490/byte_addr_base_update_enable
      -- CP-element group 5: 	 assign_stmt_322_to_assign_stmt_490/byte_addr_base_update_enable_out
      -- 
    accessMemoryByteBase_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByteBase_CP_283_elements(11);
      gj_accessMemoryByteBase_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	69 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_322_to_assign_stmt_490/offset_update_enable
      -- CP-element group 6: 	 assign_stmt_322_to_assign_stmt_490/offset_update_enable_out
      -- 
    accessMemoryByteBase_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByteBase_CP_283_elements(11);
      gj_accessMemoryByteBase_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	15 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	70 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_322_to_assign_stmt_490/wbyte_update_enable
      -- CP-element group 7: 	 assign_stmt_322_to_assign_stmt_490/wbyte_update_enable_out
      -- 
    accessMemoryByteBase_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryByteBase_CP_283_elements(15);
      gj_accessMemoryByteBase_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	71 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	62 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 assign_stmt_322_to_assign_stmt_490/rbyte_update_enable
      -- CP-element group 8: 	 assign_stmt_322_to_assign_stmt_490/rbyte_update_enable_in
      -- 
    accessMemoryByteBase_CP_283_elements(8) <= accessMemoryByteBase_CP_283_elements(71);
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_sample_start_
      -- CP-element group 9: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Sample/req
      -- 
    req_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(9), ack => call_calculateAddress36_expr_321_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "accessMemoryByteBase_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(1) & accessMemoryByteBase_CP_283_elements(11);
      gj_accessMemoryByteBase_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	27 
    -- CP-element group 10: 	31 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	39 
    -- CP-element group 10: 	43 
    -- CP-element group 10: 	47 
    -- CP-element group 10: 	51 
    -- CP-element group 10: 	55 
    -- CP-element group 10: 	59 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_update_start_
      -- CP-element group 10: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Update/$entry
      -- CP-element group 10: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Update/req
      -- 
    req_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(10), ack => call_calculateAddress36_expr_321_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(27) & accessMemoryByteBase_CP_283_elements(31) & accessMemoryByteBase_CP_283_elements(35) & accessMemoryByteBase_CP_283_elements(39) & accessMemoryByteBase_CP_283_elements(43) & accessMemoryByteBase_CP_283_elements(47) & accessMemoryByteBase_CP_283_elements(51) & accessMemoryByteBase_CP_283_elements(55) & accessMemoryByteBase_CP_283_elements(59);
      gj_accessMemoryByteBase_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_sample_completed_
      -- CP-element group 11: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Sample/ack
      -- 
    ack_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_calculateAddress36_expr_321_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	25 
    -- CP-element group 12: 	29 
    -- CP-element group 12: 	33 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	41 
    -- CP-element group 12: 	45 
    -- CP-element group 12: 	49 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	57 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_update_completed_
      -- CP-element group 12: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Update/$exit
      -- CP-element group 12: 	 assign_stmt_322_to_assign_stmt_490/call_calculateAddress36_expr_321_Update/ack
      -- 
    ack_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_calculateAddress36_expr_321_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_sample_start_
      -- CP-element group 13: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Sample/rr
      -- 
    rr_324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(13), ack => CONCAT_u8_u64_346_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(1) & accessMemoryByteBase_CP_283_elements(15);
      gj_accessMemoryByteBase_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	27 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_update_start_
      -- CP-element group 14: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Update/$entry
      -- CP-element group 14: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Update/cr
      -- 
    cr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(14), ack => CONCAT_u8_u64_346_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(16) & accessMemoryByteBase_CP_283_elements(27);
      gj_accessMemoryByteBase_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	7 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_sample_completed_
      -- CP-element group 15: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Sample/ra
      -- 
    ra_325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u64_346_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	25 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_update_completed_
      -- CP-element group 16: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Update/$exit
      -- CP-element group 16: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u8_u64_346_Update/ca
      -- 
    ca_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u64_346_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_sample_start_
      -- CP-element group 17: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Sample/rr
      -- 
    rr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(17), ack => CONCAT_u1_u2_360_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(1) & accessMemoryByteBase_CP_283_elements(19);
      gj_accessMemoryByteBase_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	27 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_update_start_
      -- CP-element group 18: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Update/$entry
      -- CP-element group 18: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Update/cr
      -- 
    cr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(18), ack => CONCAT_u1_u2_360_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(20) & accessMemoryByteBase_CP_283_elements(27);
      gj_accessMemoryByteBase_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	3 
    -- CP-element group 19: 	4 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_sample_completed_
      -- CP-element group 19: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Sample/ra
      -- 
    ra_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u2_360_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_update_completed_
      -- CP-element group 20: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Update/$exit
      -- CP-element group 20: 	 assign_stmt_322_to_assign_stmt_490/CONCAT_u1_u2_360_Update/ca
      -- 
    ca_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u2_360_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	1 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_sample_start_
      -- CP-element group 21: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Sample/req
      -- 
    req_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(21), ack => W_tag_365_delayed_3_0_371_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(1) & accessMemoryByteBase_CP_283_elements(23);
      gj_accessMemoryByteBase_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_update_start_
      -- CP-element group 22: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Update/$entry
      -- CP-element group 22: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Update/req
      -- 
    req_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(22), ack => W_tag_365_delayed_3_0_371_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(24) & accessMemoryByteBase_CP_283_elements(27);
      gj_accessMemoryByteBase_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_sample_completed_
      -- CP-element group 23: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Sample/$exit
      -- CP-element group 23: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Sample/ack
      -- 
    ack_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_365_delayed_3_0_371_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_update_completed_
      -- CP-element group 24: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Update/$exit
      -- CP-element group 24: 	 assign_stmt_322_to_assign_stmt_490/assign_stmt_373_Update/ack
      -- 
    ack_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_365_delayed_3_0_371_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	12 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	24 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_sample_start_
      -- CP-element group 25: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Sample/crr
      -- 
    crr_366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(25), ack => call_stmt_377_call_req_0); -- 
    accessMemoryByteBase_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(16) & accessMemoryByteBase_CP_283_elements(20) & accessMemoryByteBase_CP_283_elements(24) & accessMemoryByteBase_CP_283_elements(27);
      gj_accessMemoryByteBase_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: 	63 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_update_start_
      -- CP-element group 26: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Update/$entry
      -- CP-element group 26: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Update/ccr
      -- 
    ccr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(26), ack => call_stmt_377_call_req_1); -- 
    accessMemoryByteBase_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(28) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	10 
    -- CP-element group 27: 	14 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_sample_completed_
      -- CP-element group 27: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Sample/cra
      -- 
    cra_367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_377_call_ack_0, ack => accessMemoryByteBase_CP_283_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	61 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_update_completed_
      -- CP-element group 28: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Update/$exit
      -- CP-element group 28: 	 assign_stmt_322_to_assign_stmt_490/call_stmt_377_Update/cca
      -- 
    cca_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_377_call_ack_1, ack => accessMemoryByteBase_CP_283_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_sample_start_
      -- CP-element group 29: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Sample/$entry
      -- CP-element group 29: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Sample/rr
      -- 
    rr_380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(29), ack => EQ_u3_u1_413_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(31);
      gj_accessMemoryByteBase_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	63 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_update_start_
      -- CP-element group 30: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Update/$entry
      -- CP-element group 30: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Update/cr
      -- 
    cr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(30), ack => EQ_u3_u1_413_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(32) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	10 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_sample_completed_
      -- CP-element group 31: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Sample/ra
      -- 
    ra_381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_413_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	61 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_update_completed_
      -- CP-element group 32: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Update/$exit
      -- CP-element group 32: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_413_Update/ca
      -- 
    ca_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_413_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	12 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_sample_start_
      -- CP-element group 33: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Sample/$entry
      -- CP-element group 33: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Sample/rr
      -- 
    rr_394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(33), ack => EQ_u3_u1_418_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(35);
      gj_accessMemoryByteBase_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	63 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_update_start_
      -- CP-element group 34: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Update/$entry
      -- CP-element group 34: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Update/cr
      -- 
    cr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(34), ack => EQ_u3_u1_418_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(36) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_sample_completed_
      -- CP-element group 35: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Sample/ra
      -- 
    ra_395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_418_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	61 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_update_completed_
      -- CP-element group 36: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Update/$exit
      -- CP-element group 36: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_418_Update/ca
      -- 
    ca_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_418_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_sample_start_
      -- CP-element group 37: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Sample/$entry
      -- CP-element group 37: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Sample/rr
      -- 
    rr_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(37), ack => EQ_u3_u1_423_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(39);
      gj_accessMemoryByteBase_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: 	63 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_update_start_
      -- CP-element group 38: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Update/$entry
      -- CP-element group 38: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Update/cr
      -- 
    cr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(38), ack => EQ_u3_u1_423_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(40) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	10 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_sample_completed_
      -- CP-element group 39: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Sample/$exit
      -- CP-element group 39: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Sample/ra
      -- 
    ra_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_423_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	61 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_update_completed_
      -- CP-element group 40: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Update/$exit
      -- CP-element group 40: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_423_Update/ca
      -- 
    ca_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_423_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Sample/rr
      -- CP-element group 41: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Sample/$entry
      -- CP-element group 41: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_sample_start_
      -- 
    rr_422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(41), ack => EQ_u3_u1_428_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(43);
      gj_accessMemoryByteBase_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	63 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Update/$entry
      -- CP-element group 42: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Update/cr
      -- CP-element group 42: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_update_start_
      -- 
    cr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(42), ack => EQ_u3_u1_428_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(44) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	10 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Sample/ra
      -- CP-element group 43: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Sample/$exit
      -- CP-element group 43: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_sample_completed_
      -- 
    ra_423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_428_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	61 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Update/ca
      -- CP-element group 44: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_Update/$exit
      -- CP-element group 44: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_428_update_completed_
      -- 
    ca_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_428_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	12 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Sample/rr
      -- CP-element group 45: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Sample/$entry
      -- CP-element group 45: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_sample_start_
      -- 
    rr_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(45), ack => EQ_u3_u1_433_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(47);
      gj_accessMemoryByteBase_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: 	63 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Update/$entry
      -- CP-element group 46: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Update/cr
      -- CP-element group 46: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_update_start_
      -- 
    cr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(46), ack => EQ_u3_u1_433_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(48) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	10 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Sample/ra
      -- CP-element group 47: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Sample/$exit
      -- CP-element group 47: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_sample_completed_
      -- 
    ra_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_433_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(47)); -- 
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	61 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Update/$exit
      -- CP-element group 48: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_Update/ca
      -- CP-element group 48: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_433_update_completed_
      -- 
    ca_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_433_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	12 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Sample/rr
      -- CP-element group 49: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Sample/$entry
      -- CP-element group 49: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_sample_start_
      -- 
    rr_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(49), ack => EQ_u3_u1_438_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(51);
      gj_accessMemoryByteBase_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: 	63 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_update_start_
      -- CP-element group 50: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Update/cr
      -- CP-element group 50: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Update/$entry
      -- 
    cr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(50), ack => EQ_u3_u1_438_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(52) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	10 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Sample/ra
      -- CP-element group 51: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Sample/$exit
      -- CP-element group 51: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_sample_completed_
      -- 
    ra_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_438_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	61 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_update_completed_
      -- CP-element group 52: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Update/ca
      -- CP-element group 52: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_438_Update/$exit
      -- 
    ca_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_438_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Sample/$entry
      -- CP-element group 53: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_sample_start_
      -- CP-element group 53: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Sample/rr
      -- 
    rr_464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(53), ack => EQ_u3_u1_443_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(55);
      gj_accessMemoryByteBase_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	63 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_update_start_
      -- CP-element group 54: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Update/cr
      -- CP-element group 54: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Update/$entry
      -- 
    cr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(54), ack => EQ_u3_u1_443_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(56) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	10 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Sample/$exit
      -- CP-element group 55: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_sample_completed_
      -- CP-element group 55: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Sample/ra
      -- 
    ra_465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_443_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	61 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_update_completed_
      -- CP-element group 56: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Update/ca
      -- CP-element group 56: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_443_Update/$exit
      -- 
    ca_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_443_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Sample/rr
      -- CP-element group 57: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Sample/$entry
      -- CP-element group 57: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_sample_start_
      -- 
    rr_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(57), ack => EQ_u3_u1_448_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(12) & accessMemoryByteBase_CP_283_elements(59);
      gj_accessMemoryByteBase_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	63 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_update_start_
      -- CP-element group 58: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Update/cr
      -- CP-element group 58: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Update/$entry
      -- 
    cr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(58), ack => EQ_u3_u1_448_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(60) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	10 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Sample/ra
      -- CP-element group 59: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Sample/$exit
      -- CP-element group 59: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_sample_completed_
      -- 
    ra_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_448_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_update_completed_
      -- CP-element group 60: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Update/ca
      -- CP-element group 60: 	 assign_stmt_322_to_assign_stmt_490/EQ_u3_u1_448_Update/$exit
      -- 
    ca_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_448_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	28 
    -- CP-element group 61: 	32 
    -- CP-element group 61: 	36 
    -- CP-element group 61: 	40 
    -- CP-element group 61: 	44 
    -- CP-element group 61: 	48 
    -- CP-element group 61: 	52 
    -- CP-element group 61: 	56 
    -- CP-element group 61: 	60 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Sample/rr
      -- CP-element group 61: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Sample/$entry
      -- CP-element group 61: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_sample_start_
      -- 
    rr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(61), ack => OR_u8_u8_489_inst_req_0); -- 
    accessMemoryByteBase_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(28) & accessMemoryByteBase_CP_283_elements(32) & accessMemoryByteBase_CP_283_elements(36) & accessMemoryByteBase_CP_283_elements(40) & accessMemoryByteBase_CP_283_elements(44) & accessMemoryByteBase_CP_283_elements(48) & accessMemoryByteBase_CP_283_elements(52) & accessMemoryByteBase_CP_283_elements(56) & accessMemoryByteBase_CP_283_elements(60) & accessMemoryByteBase_CP_283_elements(63);
      gj_accessMemoryByteBase_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	8 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Update/cr
      -- CP-element group 62: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Update/$entry
      -- CP-element group 62: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_update_start_
      -- 
    cr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryByteBase_CP_283_elements(62), ack => OR_u8_u8_489_inst_req_1); -- 
    accessMemoryByteBase_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryByteBase_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryByteBase_CP_283_elements(8) & accessMemoryByteBase_CP_283_elements(64);
      gj_accessMemoryByteBase_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryByteBase_CP_283_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	26 
    -- CP-element group 63: 	30 
    -- CP-element group 63: 	34 
    -- CP-element group 63: 	38 
    -- CP-element group 63: 	42 
    -- CP-element group 63: 	46 
    -- CP-element group 63: 	50 
    -- CP-element group 63: 	54 
    -- CP-element group 63: 	58 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Sample/ra
      -- CP-element group 63: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Sample/$exit
      -- CP-element group 63: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_sample_completed_
      -- 
    ra_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u8_u8_489_inst_ack_0, ack => accessMemoryByteBase_CP_283_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	72 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Update/$exit
      -- CP-element group 64: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_update_completed_
      -- CP-element group 64: 	 assign_stmt_322_to_assign_stmt_490/OR_u8_u8_489_Update/ca
      -- CP-element group 64: 	 assign_stmt_322_to_assign_stmt_490/$exit
      -- 
    ca_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u8_u8_489_inst_ack_1, ack => accessMemoryByteBase_CP_283_elements(64)); -- 
    -- CP-element group 65:  place  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	2 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 tag_update_enable
      -- 
    accessMemoryByteBase_CP_283_elements(65) <= accessMemoryByteBase_CP_283_elements(2);
    -- CP-element group 66:  place  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 lock_update_enable
      -- 
    accessMemoryByteBase_CP_283_elements(66) <= accessMemoryByteBase_CP_283_elements(3);
    -- CP-element group 67:  place  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	4 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 rwbar_update_enable
      -- 
    accessMemoryByteBase_CP_283_elements(67) <= accessMemoryByteBase_CP_283_elements(4);
    -- CP-element group 68:  place  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	5 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 byte_addr_base_update_enable
      -- 
    accessMemoryByteBase_CP_283_elements(68) <= accessMemoryByteBase_CP_283_elements(5);
    -- CP-element group 69:  place  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	6 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 offset_update_enable
      -- 
    accessMemoryByteBase_CP_283_elements(69) <= accessMemoryByteBase_CP_283_elements(6);
    -- CP-element group 70:  place  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	7 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 wbyte_update_enable
      -- 
    accessMemoryByteBase_CP_283_elements(70) <= accessMemoryByteBase_CP_283_elements(7);
    -- CP-element group 71:  place  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	8 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 rbyte_update_enable
      -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	64 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 $exit
      -- 
    accessMemoryByteBase_CP_283_elements(72) <= accessMemoryByteBase_CP_283_elements(64);
    --  hookup: inputs to control-path 
    accessMemoryByteBase_CP_283_elements(71) <= rbyte_update_enable;
    -- hookup: output from control-path 
    rwbar_update_enable <= accessMemoryByteBase_CP_283_elements(67);
    lock_update_enable <= accessMemoryByteBase_CP_283_elements(66);
    offset_update_enable <= accessMemoryByteBase_CP_283_elements(69);
    byte_addr_base_update_enable <= accessMemoryByteBase_CP_283_elements(68);
    tag_update_enable <= accessMemoryByteBase_CP_283_elements(65);
    wbyte_update_enable <= accessMemoryByteBase_CP_283_elements(70);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_357_357_delayed_3_0_361 : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_365_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_368_wire : std_logic_vector(99 downto 0);
    signal CONCAT_u3_u6_353_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u8_u64_346_346_delayed_3_0_347 : std_logic_vector(63 downto 0);
    signal EQ_u3_u1_408_408_delayed_11_0_419 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_414_414_delayed_11_0_424 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_421_421_delayed_11_0_429 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_427_427_delayed_11_0_414 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_435_435_delayed_11_0_434 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_441_441_delayed_11_0_439 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_448_448_delayed_11_0_444 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_454_454_delayed_11_0_449 : std_logic_vector(0 downto 0);
    signal MUX_454_wire : std_logic_vector(7 downto 0);
    signal MUX_458_wire : std_logic_vector(7 downto 0);
    signal MUX_463_wire : std_logic_vector(7 downto 0);
    signal MUX_467_wire : std_logic_vector(7 downto 0);
    signal MUX_473_wire : std_logic_vector(7 downto 0);
    signal MUX_477_wire : std_logic_vector(7 downto 0);
    signal MUX_482_wire : std_logic_vector(7 downto 0);
    signal MUX_486_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_459_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_468_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_469_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_478_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_487_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_488_wire : std_logic_vector(7 downto 0);
    signal addr_dw_333 : std_logic_vector(35 downto 0);
    signal b0_381 : std_logic_vector(7 downto 0);
    signal b1_385 : std_logic_vector(7 downto 0);
    signal b2_389 : std_logic_vector(7 downto 0);
    signal b3_393 : std_logic_vector(7 downto 0);
    signal b4_397 : std_logic_vector(7 downto 0);
    signal b5_401 : std_logic_vector(7 downto 0);
    signal b6_405 : std_logic_vector(7 downto 0);
    signal b7_409 : std_logic_vector(7 downto 0);
    signal bb_326 : std_logic_vector(2 downto 0);
    signal bmask_340 : std_logic_vector(7 downto 0);
    signal byte_addr_322 : std_logic_vector(35 downto 0);
    signal konst_335_wire_constant : std_logic_vector(7 downto 0);
    signal konst_412_wire_constant : std_logic_vector(2 downto 0);
    signal konst_417_wire_constant : std_logic_vector(2 downto 0);
    signal konst_422_wire_constant : std_logic_vector(2 downto 0);
    signal konst_427_wire_constant : std_logic_vector(2 downto 0);
    signal konst_432_wire_constant : std_logic_vector(2 downto 0);
    signal konst_437_wire_constant : std_logic_vector(2 downto 0);
    signal konst_442_wire_constant : std_logic_vector(2 downto 0);
    signal konst_447_wire_constant : std_logic_vector(2 downto 0);
    signal konst_453_wire_constant : std_logic_vector(7 downto 0);
    signal konst_457_wire_constant : std_logic_vector(7 downto 0);
    signal konst_462_wire_constant : std_logic_vector(7 downto 0);
    signal konst_466_wire_constant : std_logic_vector(7 downto 0);
    signal konst_472_wire_constant : std_logic_vector(7 downto 0);
    signal konst_476_wire_constant : std_logic_vector(7 downto 0);
    signal konst_481_wire_constant : std_logic_vector(7 downto 0);
    signal konst_485_wire_constant : std_logic_vector(7 downto 0);
    signal request_370 : std_logic_vector(109 downto 0);
    signal response_377 : std_logic_vector(64 downto 0);
    signal slice_329_wire : std_logic_vector(32 downto 0);
    signal slice_337_wire : std_logic_vector(2 downto 0);
    signal tag_365_delayed_3_0_373 : std_logic_vector(7 downto 0);
    signal type_cast_331_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_338_wire : std_logic_vector(7 downto 0);
    signal type_cast_345_wire_constant : std_logic_vector(55 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_354_wire : std_logic_vector(63 downto 0);
    signal wdata_356 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_335_wire_constant <= "10000000";
    konst_412_wire_constant <= "011";
    konst_417_wire_constant <= "000";
    konst_422_wire_constant <= "001";
    konst_427_wire_constant <= "010";
    konst_432_wire_constant <= "100";
    konst_437_wire_constant <= "101";
    konst_442_wire_constant <= "110";
    konst_447_wire_constant <= "111";
    konst_453_wire_constant <= "00000000";
    konst_457_wire_constant <= "00000000";
    konst_462_wire_constant <= "00000000";
    konst_466_wire_constant <= "00000000";
    konst_472_wire_constant <= "00000000";
    konst_476_wire_constant <= "00000000";
    konst_481_wire_constant <= "00000000";
    konst_485_wire_constant <= "00000000";
    type_cast_331_wire_constant <= "000";
    type_cast_345_wire_constant <= "00000000000000000000000000000000000000000000000000000000";
    type_cast_352_wire_constant <= "000";
    -- flow-through select operator MUX_454_inst
    MUX_454_wire <= b0_381 when (EQ_u3_u1_408_408_delayed_11_0_419(0) /=  '0') else konst_453_wire_constant;
    -- flow-through select operator MUX_458_inst
    MUX_458_wire <= b1_385 when (EQ_u3_u1_414_414_delayed_11_0_424(0) /=  '0') else konst_457_wire_constant;
    -- flow-through select operator MUX_463_inst
    MUX_463_wire <= b2_389 when (EQ_u3_u1_421_421_delayed_11_0_429(0) /=  '0') else konst_462_wire_constant;
    -- flow-through select operator MUX_467_inst
    MUX_467_wire <= b3_393 when (EQ_u3_u1_427_427_delayed_11_0_414(0) /=  '0') else konst_466_wire_constant;
    -- flow-through select operator MUX_473_inst
    MUX_473_wire <= b4_397 when (EQ_u3_u1_435_435_delayed_11_0_434(0) /=  '0') else konst_472_wire_constant;
    -- flow-through select operator MUX_477_inst
    MUX_477_wire <= b5_401 when (EQ_u3_u1_441_441_delayed_11_0_439(0) /=  '0') else konst_476_wire_constant;
    -- flow-through select operator MUX_482_inst
    MUX_482_wire <= b6_405 when (EQ_u3_u1_448_448_delayed_11_0_444(0) /=  '0') else konst_481_wire_constant;
    -- flow-through select operator MUX_486_inst
    MUX_486_wire <= b7_409 when (EQ_u3_u1_454_454_delayed_11_0_449(0) /=  '0') else konst_485_wire_constant;
    -- flow-through slice operator slice_325_inst
    bb_326 <= byte_addr_322(2 downto 0);
    -- flow-through slice operator slice_329_inst
    slice_329_wire <= byte_addr_322(35 downto 3);
    -- flow-through slice operator slice_337_inst
    slice_337_wire <= byte_addr_322(2 downto 0);
    -- flow-through slice operator slice_380_inst
    b0_381 <= response_377(63 downto 56);
    -- flow-through slice operator slice_384_inst
    b1_385 <= response_377(55 downto 48);
    -- flow-through slice operator slice_388_inst
    b2_389 <= response_377(47 downto 40);
    -- flow-through slice operator slice_392_inst
    b3_393 <= response_377(39 downto 32);
    -- flow-through slice operator slice_396_inst
    b4_397 <= response_377(31 downto 24);
    -- flow-through slice operator slice_400_inst
    b5_401 <= response_377(23 downto 16);
    -- flow-through slice operator slice_404_inst
    b6_405 <= response_377(15 downto 8);
    -- flow-through slice operator slice_408_inst
    b7_409 <= response_377(7 downto 0);
    W_tag_365_delayed_3_0_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_tag_365_delayed_3_0_371_inst_req_0;
      W_tag_365_delayed_3_0_371_inst_ack_0<= wack(0);
      rreq(0) <= W_tag_365_delayed_3_0_371_inst_req_1;
      W_tag_365_delayed_3_0_371_inst_ack_1<= rack(0);
      W_tag_365_delayed_3_0_371_inst : InterlockBuffer generic map ( -- 
        name => "W_tag_365_delayed_3_0_371_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_365_delayed_3_0_373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_338_inst
    process(slice_337_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := slice_337_wire(2 downto 0);
      type_cast_338_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_354_inst
    process(CONCAT_u3_u6_353_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := CONCAT_u3_u6_353_wire(5 downto 0);
      type_cast_354_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator CONCAT_u10_u110_369_inst
    process(CONCAT_u2_u10_365_wire, CONCAT_u36_u100_368_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_365_wire, CONCAT_u36_u100_368_wire, tmp_var);
      request_370 <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u1_u2_360_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= lock_buffer & rwbar_buffer;
      CONCAT_u1_u2_357_357_delayed_3_0_361 <= data_out(1 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u2_360_inst_req_0;
      CONCAT_u1_u2_360_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u2_360_inst_req_1;
      CONCAT_u1_u2_360_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 2,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 3,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- flow through binary operator CONCAT_u2_u10_365_inst
    process(CONCAT_u1_u2_357_357_delayed_3_0_361, bmask_340) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_357_357_delayed_3_0_361, bmask_340, tmp_var);
      CONCAT_u2_u10_365_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u33_u36_332_inst
    process(slice_329_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_329_wire, type_cast_331_wire_constant, tmp_var);
      addr_dw_333 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u36_u100_368_inst
    process(addr_dw_333, wdata_356) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_dw_333, wdata_356, tmp_var);
      CONCAT_u36_u100_368_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u3_u6_353_inst
    process(bb_326) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(bb_326, type_cast_352_wire_constant, tmp_var);
      CONCAT_u3_u6_353_wire <= tmp_var; --
    end process;
    -- shared split operator group (6) : CONCAT_u8_u64_346_inst 
    ApConcat_group_6: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= wbyte_buffer;
      CONCAT_u8_u64_346_346_delayed_3_0_347 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u8_u64_346_inst_req_0;
      CONCAT_u8_u64_346_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u64_346_inst_req_1;
      CONCAT_u8_u64_346_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_6_gI: SplitGuardInterface generic map(name => "ApConcat_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "00000000000000000000000000000000000000000000000000000000",
          constant_width => 56,
          buffering  => 3,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u3_u1_413_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_427_427_delayed_11_0_414 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_413_inst_req_0;
      EQ_u3_u1_413_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_413_inst_req_1;
      EQ_u3_u1_413_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "011",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : EQ_u3_u1_418_inst 
    ApIntEq_group_8: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_408_408_delayed_11_0_419 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_418_inst_req_0;
      EQ_u3_u1_418_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_418_inst_req_1;
      EQ_u3_u1_418_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_8_gI: SplitGuardInterface generic map(name => "ApIntEq_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : EQ_u3_u1_423_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_414_414_delayed_11_0_424 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_423_inst_req_0;
      EQ_u3_u1_423_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_423_inst_req_1;
      EQ_u3_u1_423_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_9_gI: SplitGuardInterface generic map(name => "ApIntEq_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "001",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : EQ_u3_u1_428_inst 
    ApIntEq_group_10: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_421_421_delayed_11_0_429 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_428_inst_req_0;
      EQ_u3_u1_428_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_428_inst_req_1;
      EQ_u3_u1_428_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_10_gI: SplitGuardInterface generic map(name => "ApIntEq_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "010",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : EQ_u3_u1_433_inst 
    ApIntEq_group_11: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_435_435_delayed_11_0_434 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_433_inst_req_0;
      EQ_u3_u1_433_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_433_inst_req_1;
      EQ_u3_u1_433_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_11_gI: SplitGuardInterface generic map(name => "ApIntEq_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : EQ_u3_u1_438_inst 
    ApIntEq_group_12: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_441_441_delayed_11_0_439 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_438_inst_req_0;
      EQ_u3_u1_438_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_438_inst_req_1;
      EQ_u3_u1_438_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_12_gI: SplitGuardInterface generic map(name => "ApIntEq_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "101",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : EQ_u3_u1_443_inst 
    ApIntEq_group_13: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_448_448_delayed_11_0_444 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_443_inst_req_0;
      EQ_u3_u1_443_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_443_inst_req_1;
      EQ_u3_u1_443_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_13_gI: SplitGuardInterface generic map(name => "ApIntEq_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "110",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : EQ_u3_u1_448_inst 
    ApIntEq_group_14: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 11);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= bb_326;
      EQ_u3_u1_454_454_delayed_11_0_449 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_448_inst_req_0;
      EQ_u3_u1_448_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_448_inst_req_1;
      EQ_u3_u1_448_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_14_gI: SplitGuardInterface generic map(name => "ApIntEq_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "111",
          constant_width => 3,
          buffering  => 11,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- flow through binary operator LSHR_u64_u64_355_inst
    process(CONCAT_u8_u64_346_346_delayed_3_0_347, type_cast_354_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(CONCAT_u8_u64_346_346_delayed_3_0_347, type_cast_354_wire, tmp_var);
      wdata_356 <= tmp_var; --
    end process;
    -- flow through binary operator LSHR_u8_u8_339_inst
    process(konst_335_wire_constant, type_cast_338_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(konst_335_wire_constant, type_cast_338_wire, tmp_var);
      bmask_340 <= tmp_var; --
    end process;
    -- flow through binary operator OR_u8_u8_459_inst
    OR_u8_u8_459_wire <= (MUX_454_wire or MUX_458_wire);
    -- flow through binary operator OR_u8_u8_468_inst
    OR_u8_u8_468_wire <= (MUX_463_wire or MUX_467_wire);
    -- flow through binary operator OR_u8_u8_469_inst
    OR_u8_u8_469_wire <= (OR_u8_u8_459_wire or OR_u8_u8_468_wire);
    -- flow through binary operator OR_u8_u8_478_inst
    OR_u8_u8_478_wire <= (MUX_473_wire or MUX_477_wire);
    -- flow through binary operator OR_u8_u8_487_inst
    OR_u8_u8_487_wire <= (MUX_482_wire or MUX_486_wire);
    -- flow through binary operator OR_u8_u8_488_inst
    OR_u8_u8_488_wire <= (OR_u8_u8_478_wire or OR_u8_u8_487_wire);
    -- shared split operator group (23) : OR_u8_u8_489_inst 
    ApIntOr_group_23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OR_u8_u8_469_wire & OR_u8_u8_488_wire;
      rbyte_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u8_u8_489_inst_req_0;
      OR_u8_u8_489_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u8_u8_489_inst_req_1;
      OR_u8_u8_489_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_23_gI: SplitGuardInterface generic map(name => "ApIntOr_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared call operator group (0) : call_calculateAddress36_expr_321_inst 
    calculateAddress36_call_group_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_calculateAddress36_expr_321_inst_req_0;
      call_calculateAddress36_expr_321_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_calculateAddress36_expr_321_inst_req_1;
      call_calculateAddress36_expr_321_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      calculateAddress36_call_group_0_gI: SplitGuardInterface generic map(name => "calculateAddress36_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= byte_addr_base_buffer & offset_buffer;
      byte_addr_322 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => calculateAddress36_call_reqs(0),
          ackR => calculateAddress36_call_acks(0),
          dataR => calculateAddress36_call_data(127 downto 0),
          tagR => calculateAddress36_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => calculateAddress36_return_acks(0), -- cross-over
          ackL => calculateAddress36_return_reqs(0), -- cross-over
          dataL => calculateAddress36_return_data(35 downto 0),
          tagL => calculateAddress36_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_377_call 
    accessMemoryBase_call_group_1: Block -- 
      signal data_in: std_logic_vector(117 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 11);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_377_call_req_0;
      call_stmt_377_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_377_call_req_1;
      call_stmt_377_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryBase_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryBase_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_365_delayed_3_0_373 & request_370;
      response_377 <= data_out(64 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 118,
        owidth => 118,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryBase_call_reqs(0),
          ackR => accessMemoryBase_call_acks(0),
          dataR => accessMemoryBase_call_data(117 downto 0),
          tagR => accessMemoryBase_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 65,
          owidth => 65,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryBase_return_acks(0), -- cross-over
          ackL => accessMemoryBase_return_reqs(0), -- cross-over
          dataL => accessMemoryBase_return_data(64 downto 0),
          tagL => accessMemoryBase_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end accessMemoryByteBase_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryDword is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    base_addr : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_call_data : out  std_logic_vector(202 downto 0);
    doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
    doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_return_data : in   std_logic_vector(63 downto 0);
    doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryDword;
architecture accessMemoryDword_arch of accessMemoryDword is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 201)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal base_addr_buffer :  std_logic_vector(63 downto 0);
  signal base_addr_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemoryDword_CP_1479_start: Boolean;
  signal accessMemoryDword_CP_1479_symbol: Boolean;
  -- volatile/operator module components. 
  component doMemAccess is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      opcode : in  std_logic_vector(2 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      memory_access_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_data : out  std_logic_vector(169 downto 0);
      accessMemoryWordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWordBase_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_data : out  std_logic_vector(145 downto 0);
      accessMemoryByteBase_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryByteBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByteBase_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemoryDwordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_data : out  std_logic_vector(201 downto 0);
      accessMemoryDwordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDwordBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1089_call_req_0 : boolean;
  signal call_stmt_1089_call_ack_0 : boolean;
  signal call_stmt_1089_call_ack_1 : boolean;
  signal call_stmt_1089_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryDword_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 201) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= base_addr;
  base_addr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(136 downto 73) <= offset;
  offset_buffer <= in_buffer_data_out(136 downto 73);
  in_buffer_data_in(200 downto 137) <= wdata;
  wdata_buffer <= in_buffer_data_out(200 downto 137);
  in_buffer_data_in(tag_length + 200 downto 201) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 200 downto 201);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 1,6 => 7);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 7);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= tag_update_enable & rwbar_update_enable & base_addr_update_enable & offset_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryDword_CP_1479_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryDword_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryDword_CP_1479_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryDword_CP_1479_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryDword_CP_1479_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryDword_CP_1479: Block -- control-path 
    signal accessMemoryDword_CP_1479_elements: BooleanArray(18 downto 0);
    -- 
  begin -- 
    accessMemoryDword_CP_1479_elements(0) <= accessMemoryDword_CP_1479_start;
    accessMemoryDword_CP_1479_symbol <= accessMemoryDword_CP_1479_elements(18);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1089/$entry
      -- 
    accessMemoryDword_CP_1479_elements(1) <= accessMemoryDword_CP_1479_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1089/tag_update_enable_out
      -- CP-element group 2: 	 call_stmt_1089/tag_update_enable
      -- 
    accessMemoryDword_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDword_CP_1479_elements(10);
      gj_accessMemoryDword_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	10 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1089/rwbar_update_enable
      -- CP-element group 3: 	 call_stmt_1089/rwbar_update_enable_out
      -- 
    accessMemoryDword_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDword_CP_1479_elements(10);
      gj_accessMemoryDword_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	10 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	14 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_1089/base_addr_update_enable_out
      -- CP-element group 4: 	 call_stmt_1089/base_addr_update_enable
      -- 
    accessMemoryDword_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDword_CP_1479_elements(10);
      gj_accessMemoryDword_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	15 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_1089/offset_update_enable_out
      -- CP-element group 5: 	 call_stmt_1089/offset_update_enable
      -- 
    accessMemoryDword_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDword_CP_1479_elements(10);
      gj_accessMemoryDword_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	10 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	16 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 call_stmt_1089/wdata_update_enable_out
      -- CP-element group 6: 	 call_stmt_1089/wdata_update_enable
      -- 
    accessMemoryDword_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDword_CP_1479_elements(10);
      gj_accessMemoryDword_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	17 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 call_stmt_1089/rdata_update_enable
      -- CP-element group 7: 	 call_stmt_1089/rdata_update_enable_in
      -- 
    accessMemoryDword_CP_1479_elements(7) <= accessMemoryDword_CP_1479_elements(17);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1089/call_stmt_1089_sample_start_
      -- CP-element group 8: 	 call_stmt_1089/call_stmt_1089_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1089/call_stmt_1089_Sample/crr
      -- 
    crr_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDword_CP_1479_elements(8), ack => call_stmt_1089_call_req_0); -- 
    accessMemoryDword_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDword_CP_1479_elements(1) & accessMemoryDword_CP_1479_elements(10);
      gj_accessMemoryDword_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1089/call_stmt_1089_Update/$entry
      -- CP-element group 9: 	 call_stmt_1089/call_stmt_1089_update_start_
      -- CP-element group 9: 	 call_stmt_1089/call_stmt_1089_Update/ccr
      -- 
    ccr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDword_CP_1479_elements(9), ack => call_stmt_1089_call_req_1); -- 
    accessMemoryDword_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "accessMemoryDword_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDword_CP_1479_elements(7) & accessMemoryDword_CP_1479_elements(11);
      gj_accessMemoryDword_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDword_CP_1479_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: 	5 
    -- CP-element group 10: 	6 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1089/call_stmt_1089_sample_completed_
      -- CP-element group 10: 	 call_stmt_1089/call_stmt_1089_Sample/$exit
      -- CP-element group 10: 	 call_stmt_1089/call_stmt_1089_Sample/cra
      -- 
    cra_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1089_call_ack_0, ack => accessMemoryDword_CP_1479_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	18 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 call_stmt_1089/call_stmt_1089_Update/$exit
      -- CP-element group 11: 	 call_stmt_1089/$exit
      -- CP-element group 11: 	 call_stmt_1089/call_stmt_1089_update_completed_
      -- CP-element group 11: 	 call_stmt_1089/call_stmt_1089_Update/cca
      -- 
    cca_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1089_call_ack_1, ack => accessMemoryDword_CP_1479_elements(11)); -- 
    -- CP-element group 12:  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 tag_update_enable
      -- 
    accessMemoryDword_CP_1479_elements(12) <= accessMemoryDword_CP_1479_elements(2);
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 rwbar_update_enable
      -- 
    accessMemoryDword_CP_1479_elements(13) <= accessMemoryDword_CP_1479_elements(3);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	4 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 base_addr_update_enable
      -- 
    accessMemoryDword_CP_1479_elements(14) <= accessMemoryDword_CP_1479_elements(4);
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	5 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 offset_update_enable
      -- 
    accessMemoryDword_CP_1479_elements(15) <= accessMemoryDword_CP_1479_elements(5);
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	6 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 wdata_update_enable
      -- 
    accessMemoryDword_CP_1479_elements(16) <= accessMemoryDword_CP_1479_elements(6);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	7 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rdata_update_enable
      -- 
    -- CP-element group 18:  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 $exit
      -- 
    accessMemoryDword_CP_1479_elements(18) <= accessMemoryDword_CP_1479_elements(11);
    --  hookup: inputs to control-path 
    accessMemoryDword_CP_1479_elements(17) <= rdata_update_enable;
    -- hookup: output from control-path 
    wdata_update_enable <= accessMemoryDword_CP_1479_elements(16);
    offset_update_enable <= accessMemoryDword_CP_1479_elements(15);
    base_addr_update_enable <= accessMemoryDword_CP_1479_elements(14);
    rwbar_update_enable <= accessMemoryDword_CP_1479_elements(13);
    tag_update_enable <= accessMemoryDword_CP_1479_elements(12);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_1084_wire : std_logic_vector(2 downto 0);
    signal R_LDD_1082_wire_constant : std_logic_vector(2 downto 0);
    signal R_STD_1083_wire_constant : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    R_LDD_1082_wire_constant <= "101";
    R_STD_1083_wire_constant <= "010";
    -- flow-through select operator MUX_1084_inst
    MUX_1084_wire <= R_LDD_1082_wire_constant when (rwbar_buffer(0) /=  '0') else R_STD_1083_wire_constant;
    -- shared call operator group (0) : call_stmt_1089_call 
    doMemAccess_call_group_0: Block -- 
      signal data_in: std_logic_vector(202 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 36);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1089_call_req_0;
      call_stmt_1089_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1089_call_req_1;
      call_stmt_1089_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      doMemAccess_call_group_0_gI: SplitGuardInterface generic map(name => "doMemAccess_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & MUX_1084_wire & base_addr_buffer & offset_buffer & wdata_buffer;
      rdata_buffer <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 203,
        owidth => 203,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => doMemAccess_call_reqs(0),
          ackR => doMemAccess_call_acks(0),
          dataR => doMemAccess_call_data(202 downto 0),
          tagR => doMemAccess_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => doMemAccess_return_acks(0), -- cross-over
          ackL => doMemAccess_return_reqs(0), -- cross-over
          dataL => doMemAccess_return_data(63 downto 0),
          tagL => doMemAccess_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemoryDword_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryDwordBase is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    base_addr : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
    calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
    calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
    calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
    calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
    calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
    calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
    calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
    accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
    accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryDwordBase;
architecture accessMemoryDwordBase_arch of accessMemoryDwordBase is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 202)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal base_addr_buffer :  std_logic_vector(63 downto 0);
  signal base_addr_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemoryDwordBase_CP_645_start: Boolean;
  signal accessMemoryDwordBase_CP_645_symbol: Boolean;
  -- volatile/operator module components. 
  component calculateAddress36 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      addr : out  std_logic_vector(35 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      request : in  std_logic_vector(109 downto 0);
      response : out  std_logic_vector(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_data : out  std_logic_vector(255 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_tag_567_delayed_3_0_613_inst_ack_1 : boolean;
  signal W_wdata_563_delayed_3_0_603_inst_req_0 : boolean;
  signal W_wdata_563_delayed_3_0_603_inst_ack_0 : boolean;
  signal W_tag_567_delayed_3_0_613_inst_req_0 : boolean;
  signal W_tag_567_delayed_3_0_613_inst_ack_0 : boolean;
  signal W_tag_567_delayed_3_0_613_inst_req_1 : boolean;
  signal call_calculateAddress36_expr_592_inst_req_1 : boolean;
  signal call_stmt_619_call_ack_0 : boolean;
  signal call_calculateAddress36_expr_592_inst_req_0 : boolean;
  signal call_calculateAddress36_expr_592_inst_ack_0 : boolean;
  signal W_wdata_563_delayed_3_0_603_inst_ack_1 : boolean;
  signal call_stmt_619_call_req_1 : boolean;
  signal call_calculateAddress36_expr_592_inst_ack_1 : boolean;
  signal call_stmt_619_call_ack_1 : boolean;
  signal W_wdata_563_delayed_3_0_603_inst_req_1 : boolean;
  signal CONCAT_u2_u10_601_inst_req_0 : boolean;
  signal call_stmt_619_call_req_0 : boolean;
  signal CONCAT_u2_u10_601_inst_ack_1 : boolean;
  signal CONCAT_u2_u10_601_inst_req_1 : boolean;
  signal CONCAT_u2_u10_601_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryDwordBase_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 202) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= lock;
  lock_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(9 downto 9) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(9 downto 9);
  in_buffer_data_in(73 downto 10) <= base_addr;
  base_addr_buffer <= in_buffer_data_out(73 downto 10);
  in_buffer_data_in(137 downto 74) <= offset;
  offset_buffer <= in_buffer_data_out(137 downto 74);
  in_buffer_data_in(201 downto 138) <= wdata;
  wdata_buffer <= in_buffer_data_out(201 downto 138);
  in_buffer_data_in(tag_length + 201 downto 202) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 201 downto 202);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 1,7 => 7);
    constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1,7 => 7);
    constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 8); -- 
  begin -- 
    preds <= tag_update_enable & lock_update_enable & rwbar_update_enable & base_addr_update_enable & offset_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryDwordBase_CP_645_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryDwordBase_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryDwordBase_CP_645_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryDwordBase_CP_645_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryDwordBase_CP_645_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryDwordBase_CP_645: Block -- control-path 
    signal accessMemoryDwordBase_CP_645_elements: BooleanArray(36 downto 0);
    -- 
  begin -- 
    accessMemoryDwordBase_CP_645_elements(0) <= accessMemoryDwordBase_CP_645_start;
    accessMemoryDwordBase_CP_645_symbol <= accessMemoryDwordBase_CP_645_elements(36);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	21 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_593_to_assign_stmt_623/$entry
      -- 
    accessMemoryDwordBase_CP_645_elements(1) <= accessMemoryDwordBase_CP_645_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	23 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	29 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_593_to_assign_stmt_623/tag_update_enable
      -- CP-element group 2: 	 assign_stmt_593_to_assign_stmt_623/tag_update_enable_out
      -- 
    accessMemoryDwordBase_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDwordBase_CP_645_elements(23);
      gj_accessMemoryDwordBase_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	30 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_593_to_assign_stmt_623/lock_update_enable_out
      -- CP-element group 3: 	 assign_stmt_593_to_assign_stmt_623/lock_update_enable
      -- 
    accessMemoryDwordBase_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDwordBase_CP_645_elements(15);
      gj_accessMemoryDwordBase_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	31 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_593_to_assign_stmt_623/rwbar_update_enable
      -- CP-element group 4: 	 assign_stmt_593_to_assign_stmt_623/rwbar_update_enable_out
      -- 
    accessMemoryDwordBase_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDwordBase_CP_645_elements(15);
      gj_accessMemoryDwordBase_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	32 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_593_to_assign_stmt_623/base_addr_update_enable
      -- CP-element group 5: 	 assign_stmt_593_to_assign_stmt_623/base_addr_update_enable_out
      -- 
    accessMemoryDwordBase_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDwordBase_CP_645_elements(11);
      gj_accessMemoryDwordBase_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	33 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_593_to_assign_stmt_623/offset_update_enable
      -- CP-element group 6: 	 assign_stmt_593_to_assign_stmt_623/offset_update_enable_out
      -- 
    accessMemoryDwordBase_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDwordBase_CP_645_elements(11);
      gj_accessMemoryDwordBase_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	34 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_593_to_assign_stmt_623/wdata_update_enable
      -- CP-element group 7: 	 assign_stmt_593_to_assign_stmt_623/wdata_update_enable_out
      -- 
    accessMemoryDwordBase_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryDwordBase_CP_645_elements(19);
      gj_accessMemoryDwordBase_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	35 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	26 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 assign_stmt_593_to_assign_stmt_623/rdata_update_enable_in
      -- CP-element group 8: 	 assign_stmt_593_to_assign_stmt_623/rdata_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(8) <= accessMemoryDwordBase_CP_645_elements(35);
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Sample/req
      -- CP-element group 9: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_sample_start_
      -- CP-element group 9: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Sample/$entry
      -- 
    req_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(9), ack => call_calculateAddress36_expr_592_inst_req_0); -- 
    accessMemoryDwordBase_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryDwordBase_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(1) & accessMemoryDwordBase_CP_645_elements(11);
      gj_accessMemoryDwordBase_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	27 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Update/req
      -- CP-element group 10: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Update/$entry
      -- CP-element group 10: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_update_start_
      -- 
    req_677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(10), ack => call_calculateAddress36_expr_592_inst_req_1); -- 
    accessMemoryDwordBase_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(12) & accessMemoryDwordBase_CP_645_elements(27);
      gj_accessMemoryDwordBase_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Sample/ack
      -- CP-element group 11: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_sample_completed_
      -- 
    ack_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_calculateAddress36_expr_592_inst_ack_0, ack => accessMemoryDwordBase_CP_645_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	25 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Update/$exit
      -- CP-element group 12: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_Update/ack
      -- CP-element group 12: 	 assign_stmt_593_to_assign_stmt_623/call_calculateAddress36_expr_592_update_completed_
      -- 
    ack_678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_calculateAddress36_expr_592_inst_ack_1, ack => accessMemoryDwordBase_CP_645_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_sample_start_
      -- CP-element group 13: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Sample/rr
      -- 
    rr_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(13), ack => CONCAT_u2_u10_601_inst_req_0); -- 
    accessMemoryDwordBase_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(1) & accessMemoryDwordBase_CP_645_elements(15);
      gj_accessMemoryDwordBase_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	27 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_update_start_
      -- CP-element group 14: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Update/cr
      -- CP-element group 14: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Update/$entry
      -- 
    cr_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(14), ack => CONCAT_u2_u10_601_inst_req_1); -- 
    accessMemoryDwordBase_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(16) & accessMemoryDwordBase_CP_645_elements(27);
      gj_accessMemoryDwordBase_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	3 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_sample_completed_
      -- CP-element group 15: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Sample/ra
      -- 
    ra_687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u2_u10_601_inst_ack_0, ack => accessMemoryDwordBase_CP_645_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	25 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_update_completed_
      -- CP-element group 16: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Update/ca
      -- CP-element group 16: 	 assign_stmt_593_to_assign_stmt_623/CONCAT_u2_u10_601_Update/$exit
      -- 
    ca_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u2_u10_601_inst_ack_1, ack => accessMemoryDwordBase_CP_645_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Sample/req
      -- CP-element group 17: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_sample_start_
      -- 
    req_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(17), ack => W_wdata_563_delayed_3_0_603_inst_req_0); -- 
    accessMemoryDwordBase_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(1) & accessMemoryDwordBase_CP_645_elements(19);
      gj_accessMemoryDwordBase_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	27 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Update/$entry
      -- CP-element group 18: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Update/req
      -- CP-element group 18: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_update_start_
      -- 
    req_705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(18), ack => W_wdata_563_delayed_3_0_603_inst_req_1); -- 
    accessMemoryDwordBase_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(20) & accessMemoryDwordBase_CP_645_elements(27);
      gj_accessMemoryDwordBase_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Sample/ack
      -- CP-element group 19: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_sample_completed_
      -- 
    ack_701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_563_delayed_3_0_603_inst_ack_0, ack => accessMemoryDwordBase_CP_645_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Update/$exit
      -- CP-element group 20: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_Update/ack
      -- CP-element group 20: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_605_update_completed_
      -- 
    ack_706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_563_delayed_3_0_603_inst_ack_1, ack => accessMemoryDwordBase_CP_645_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	1 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Sample/req
      -- CP-element group 21: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_sample_start_
      -- 
    req_714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(21), ack => W_tag_567_delayed_3_0_613_inst_req_0); -- 
    accessMemoryDwordBase_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(1) & accessMemoryDwordBase_CP_645_elements(23);
      gj_accessMemoryDwordBase_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Update/req
      -- CP-element group 22: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Update/$entry
      -- CP-element group 22: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_update_start_
      -- 
    req_719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(22), ack => W_tag_567_delayed_3_0_613_inst_req_1); -- 
    accessMemoryDwordBase_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(24) & accessMemoryDwordBase_CP_645_elements(27);
      gj_accessMemoryDwordBase_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Sample/ack
      -- CP-element group 23: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_sample_completed_
      -- CP-element group 23: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Sample/$exit
      -- 
    ack_715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_567_delayed_3_0_613_inst_ack_0, ack => accessMemoryDwordBase_CP_645_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Update/ack
      -- CP-element group 24: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_update_completed_
      -- CP-element group 24: 	 assign_stmt_593_to_assign_stmt_623/assign_stmt_615_Update/$exit
      -- 
    ack_720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_567_delayed_3_0_613_inst_ack_1, ack => accessMemoryDwordBase_CP_645_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	12 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	24 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_sample_start_
      -- CP-element group 25: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Sample/crr
      -- 
    crr_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(25), ack => call_stmt_619_call_req_0); -- 
    accessMemoryDwordBase_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(12) & accessMemoryDwordBase_CP_645_elements(16) & accessMemoryDwordBase_CP_645_elements(20) & accessMemoryDwordBase_CP_645_elements(24) & accessMemoryDwordBase_CP_645_elements(27);
      gj_accessMemoryDwordBase_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	8 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Update/$entry
      -- CP-element group 26: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Update/ccr
      -- CP-element group 26: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_update_start_
      -- 
    ccr_733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryDwordBase_CP_645_elements(26), ack => call_stmt_619_call_req_1); -- 
    accessMemoryDwordBase_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 41) := "accessMemoryDwordBase_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryDwordBase_CP_645_elements(8) & accessMemoryDwordBase_CP_645_elements(28);
      gj_accessMemoryDwordBase_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryDwordBase_CP_645_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	10 
    -- CP-element group 27: 	14 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Sample/cra
      -- CP-element group 27: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_sample_completed_
      -- CP-element group 27: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Sample/$exit
      -- 
    cra_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_619_call_ack_0, ack => accessMemoryDwordBase_CP_645_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	36 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 assign_stmt_593_to_assign_stmt_623/$exit
      -- CP-element group 28: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Update/cca
      -- CP-element group 28: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_Update/$exit
      -- CP-element group 28: 	 assign_stmt_593_to_assign_stmt_623/call_stmt_619_update_completed_
      -- 
    cca_734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_619_call_ack_1, ack => accessMemoryDwordBase_CP_645_elements(28)); -- 
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 tag_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(29) <= accessMemoryDwordBase_CP_645_elements(2);
    -- CP-element group 30:  place  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	3 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 lock_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(30) <= accessMemoryDwordBase_CP_645_elements(3);
    -- CP-element group 31:  place  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	4 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 rwbar_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(31) <= accessMemoryDwordBase_CP_645_elements(4);
    -- CP-element group 32:  place  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	5 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 base_addr_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(32) <= accessMemoryDwordBase_CP_645_elements(5);
    -- CP-element group 33:  place  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	6 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 offset_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(33) <= accessMemoryDwordBase_CP_645_elements(6);
    -- CP-element group 34:  place  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	7 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 wdata_update_enable
      -- 
    accessMemoryDwordBase_CP_645_elements(34) <= accessMemoryDwordBase_CP_645_elements(7);
    -- CP-element group 35:  place  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	8 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 rdata_update_enable
      -- 
    -- CP-element group 36:  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	28 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 $exit
      -- 
    accessMemoryDwordBase_CP_645_elements(36) <= accessMemoryDwordBase_CP_645_elements(28);
    --  hookup: inputs to control-path 
    accessMemoryDwordBase_CP_645_elements(35) <= rdata_update_enable;
    -- hookup: output from control-path 
    wdata_update_enable <= accessMemoryDwordBase_CP_645_elements(34);
    base_addr_update_enable <= accessMemoryDwordBase_CP_645_elements(32);
    offset_update_enable <= accessMemoryDwordBase_CP_645_elements(33);
    rwbar_update_enable <= accessMemoryDwordBase_CP_645_elements(31);
    lock_update_enable <= accessMemoryDwordBase_CP_645_elements(30);
    tag_update_enable <= accessMemoryDwordBase_CP_645_elements(29);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_597_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_561_561_delayed_3_0_602 : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_610_wire : std_logic_vector(99 downto 0);
    signal NOT_u8_u8_600_wire_constant : std_logic_vector(7 downto 0);
    signal addr_593 : std_logic_vector(35 downto 0);
    signal request_612 : std_logic_vector(109 downto 0);
    signal response_619 : std_logic_vector(64 downto 0);
    signal tag_567_delayed_3_0_615 : std_logic_vector(7 downto 0);
    signal wdata_563_delayed_3_0_605 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_600_wire_constant <= "11111111";
    -- flow-through slice operator slice_622_inst
    rdata_buffer <= response_619(63 downto 0);
    W_tag_567_delayed_3_0_613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_tag_567_delayed_3_0_613_inst_req_0;
      W_tag_567_delayed_3_0_613_inst_ack_0<= wack(0);
      rreq(0) <= W_tag_567_delayed_3_0_613_inst_req_1;
      W_tag_567_delayed_3_0_613_inst_ack_1<= rack(0);
      W_tag_567_delayed_3_0_613_inst : InterlockBuffer generic map ( -- 
        name => "W_tag_567_delayed_3_0_613_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_567_delayed_3_0_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_563_delayed_3_0_603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_563_delayed_3_0_603_inst_req_0;
      W_wdata_563_delayed_3_0_603_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_563_delayed_3_0_603_inst_req_1;
      W_wdata_563_delayed_3_0_603_inst_ack_1<= rack(0);
      W_wdata_563_delayed_3_0_603_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_563_delayed_3_0_603_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_563_delayed_3_0_605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- flow through binary operator CONCAT_u10_u110_611_inst
    process(CONCAT_u2_u10_561_561_delayed_3_0_602, CONCAT_u36_u100_610_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_561_561_delayed_3_0_602, CONCAT_u36_u100_610_wire, tmp_var);
      request_612 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u2_597_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_597_wire <= tmp_var; --
    end process;
    -- shared split operator group (2) : CONCAT_u2_u10_601_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(9 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u2_597_wire;
      CONCAT_u2_u10_561_561_delayed_3_0_602 <= data_out(9 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u2_u10_601_inst_req_0;
      CONCAT_u2_u10_601_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u2_u10_601_inst_req_1;
      CONCAT_u2_u10_601_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 10,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 3,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- flow through binary operator CONCAT_u36_u100_610_inst
    process(addr_593, wdata_563_delayed_3_0_605) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_593, wdata_563_delayed_3_0_605, tmp_var);
      CONCAT_u36_u100_610_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_calculateAddress36_expr_592_inst 
    calculateAddress36_call_group_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_calculateAddress36_expr_592_inst_req_0;
      call_calculateAddress36_expr_592_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_calculateAddress36_expr_592_inst_req_1;
      call_calculateAddress36_expr_592_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      calculateAddress36_call_group_0_gI: SplitGuardInterface generic map(name => "calculateAddress36_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= base_addr_buffer & offset_buffer;
      addr_593 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => calculateAddress36_call_reqs(0),
          ackR => calculateAddress36_call_acks(0),
          dataR => calculateAddress36_call_data(127 downto 0),
          tagR => calculateAddress36_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => calculateAddress36_return_acks(0), -- cross-over
          ackL => calculateAddress36_return_reqs(0), -- cross-over
          dataL => calculateAddress36_return_data(35 downto 0),
          tagL => calculateAddress36_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_619_call 
    accessMemoryBase_call_group_1: Block -- 
      signal data_in: std_logic_vector(117 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 11);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_619_call_req_0;
      call_stmt_619_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_619_call_req_1;
      call_stmt_619_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryBase_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryBase_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_567_delayed_3_0_615 & request_612;
      response_619 <= data_out(64 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 118,
        owidth => 118,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryBase_call_reqs(0),
          ackR => accessMemoryBase_call_acks(0),
          dataR => accessMemoryBase_call_data(117 downto 0),
          tagR => accessMemoryBase_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 65,
          owidth => 65,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryBase_return_acks(0), -- cross-over
          ackL => accessMemoryBase_return_reqs(0), -- cross-over
          dataL => accessMemoryBase_return_data(64 downto 0),
          tagL => accessMemoryBase_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end accessMemoryDwordBase_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryLdStub is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    byte_addr_base : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    rbyte : out  std_logic_vector(7 downto 0);
    doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_call_data : out  std_logic_vector(202 downto 0);
    doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
    doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_return_data : in   std_logic_vector(63 downto 0);
    doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryLdStub;
architecture accessMemoryLdStub_arch of accessMemoryLdStub is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 136)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal byte_addr_base_buffer :  std_logic_vector(63 downto 0);
  signal byte_addr_base_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  -- output port buffer signals
  signal rbyte_buffer :  std_logic_vector(7 downto 0);
  signal rbyte_update_enable: Boolean;
  signal accessMemoryLdStub_CP_1142_start: Boolean;
  signal accessMemoryLdStub_CP_1142_symbol: Boolean;
  -- volatile/operator module components. 
  component doMemAccess is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      opcode : in  std_logic_vector(2 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      memory_access_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_data : out  std_logic_vector(169 downto 0);
      accessMemoryWordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWordBase_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_data : out  std_logic_vector(145 downto 0);
      accessMemoryByteBase_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryByteBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByteBase_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemoryDwordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_data : out  std_logic_vector(201 downto 0);
      accessMemoryDwordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDwordBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal slice_914_inst_req_1 : boolean;
  signal call_stmt_911_call_ack_0 : boolean;
  signal call_stmt_911_call_req_1 : boolean;
  signal slice_914_inst_ack_1 : boolean;
  signal call_stmt_911_call_req_0 : boolean;
  signal slice_914_inst_ack_0 : boolean;
  signal call_stmt_911_call_ack_1 : boolean;
  signal slice_914_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryLdStub_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 136) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= byte_addr_base;
  byte_addr_base_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(135 downto 72) <= offset;
  offset_buffer <= in_buffer_data_out(135 downto 72);
  in_buffer_data_in(tag_length + 135 downto 136) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 135 downto 136);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryLdStub_CP_1142_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryLdStub_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= rbyte_buffer;
  rbyte <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryLdStub_CP_1142_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryLdStub_CP_1142_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryLdStub_CP_1142_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryLdStub_CP_1142: Block -- control-path 
    signal accessMemoryLdStub_CP_1142_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    accessMemoryLdStub_CP_1142_elements(0) <= accessMemoryLdStub_CP_1142_start;
    accessMemoryLdStub_CP_1142_symbol <= accessMemoryLdStub_CP_1142_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/slice_914_Update/cr
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Update/$entry
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_update_start_
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_sample_start_
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/$entry
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/slice_914_Update/$entry
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Sample/$entry
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Sample/crr
      -- CP-element group 0: 	 call_stmt_911_to_assign_stmt_915/slice_914_update_start_
      -- 
    crr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryLdStub_CP_1142_elements(0), ack => call_stmt_911_call_req_0); -- 
    ccr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryLdStub_CP_1142_elements(0), ack => call_stmt_911_call_req_1); -- 
    cr_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryLdStub_CP_1142_elements(0), ack => slice_914_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Sample/cra
      -- CP-element group 1: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_sample_completed_
      -- CP-element group 1: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Sample/$exit
      -- 
    cra_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_911_call_ack_0, ack => accessMemoryLdStub_CP_1142_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_update_completed_
      -- CP-element group 2: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Update/$exit
      -- CP-element group 2: 	 call_stmt_911_to_assign_stmt_915/slice_914_sample_start_
      -- CP-element group 2: 	 call_stmt_911_to_assign_stmt_915/call_stmt_911_Update/cca
      -- CP-element group 2: 	 call_stmt_911_to_assign_stmt_915/slice_914_Sample/rr
      -- CP-element group 2: 	 call_stmt_911_to_assign_stmt_915/slice_914_Sample/$entry
      -- 
    cca_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_911_call_ack_1, ack => accessMemoryLdStub_CP_1142_elements(2)); -- 
    rr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryLdStub_CP_1142_elements(2), ack => slice_914_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_911_to_assign_stmt_915/slice_914_Sample/ra
      -- CP-element group 3: 	 call_stmt_911_to_assign_stmt_915/slice_914_sample_completed_
      -- CP-element group 3: 	 call_stmt_911_to_assign_stmt_915/slice_914_Sample/$exit
      -- 
    ra_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_914_inst_ack_0, ack => accessMemoryLdStub_CP_1142_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 call_stmt_911_to_assign_stmt_915/$exit
      -- CP-element group 4: 	 call_stmt_911_to_assign_stmt_915/slice_914_Update/$exit
      -- CP-element group 4: 	 call_stmt_911_to_assign_stmt_915/slice_914_Update/ca
      -- CP-element group 4: 	 call_stmt_911_to_assign_stmt_915/slice_914_update_completed_
      -- CP-element group 4: 	 $exit
      -- 
    ca_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_914_inst_ack_1, ack => accessMemoryLdStub_CP_1142_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_LDSTUB_905_wire_constant : std_logic_vector(2 downto 0);
    signal rdword_911 : std_logic_vector(63 downto 0);
    signal type_cast_909_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    R_LDSTUB_905_wire_constant <= "111";
    type_cast_909_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_914_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_914_inst_req_0;
      slice_914_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_914_inst_req_1;
      slice_914_inst_ack_1<= update_ack(0);
      slice_914_inst: SliceSplitProtocol generic map(name => "slice_914_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdword_911, dout => rbyte_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared call operator group (0) : call_stmt_911_call 
    doMemAccess_call_group_0: Block -- 
      signal data_in: std_logic_vector(202 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_911_call_req_0;
      call_stmt_911_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_911_call_req_1;
      call_stmt_911_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      doMemAccess_call_group_0_gI: SplitGuardInterface generic map(name => "doMemAccess_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_LDSTUB_905_wire_constant & byte_addr_base_buffer & offset_buffer & type_cast_909_wire_constant;
      rdword_911 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 203,
        owidth => 203,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => doMemAccess_call_reqs(0),
          ackR => doMemAccess_call_acks(0),
          dataR => doMemAccess_call_data(202 downto 0),
          tagR => doMemAccess_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => doMemAccess_return_acks(0), -- cross-over
          ackL => doMemAccess_return_reqs(0), -- cross-over
          dataL => doMemAccess_return_data(63 downto 0),
          tagL => doMemAccess_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemoryLdStub_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryWord is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    word_addr_base : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wword : in  std_logic_vector(31 downto 0);
    rword : out  std_logic_vector(31 downto 0);
    doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_call_data : out  std_logic_vector(202 downto 0);
    doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
    doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
    doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
    doMemAccess_return_data : in   std_logic_vector(63 downto 0);
    doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryWord;
architecture accessMemoryWord_arch of accessMemoryWord is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 169)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal word_addr_base_buffer :  std_logic_vector(63 downto 0);
  signal word_addr_base_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wword_buffer :  std_logic_vector(31 downto 0);
  signal wword_update_enable: Boolean;
  -- output port buffer signals
  signal rword_buffer :  std_logic_vector(31 downto 0);
  signal rword_update_enable: Boolean;
  signal accessMemoryWord_CP_1007_start: Boolean;
  signal accessMemoryWord_CP_1007_symbol: Boolean;
  -- volatile/operator module components. 
  component doMemAccess is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      opcode : in  std_logic_vector(2 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      memory_access_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_data : out  std_logic_vector(169 downto 0);
      accessMemoryWordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWordBase_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_data : out  std_logic_vector(145 downto 0);
      accessMemoryByteBase_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryByteBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByteBase_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemoryDwordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_data : out  std_logic_vector(201 downto 0);
      accessMemoryDwordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDwordBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_846_call_ack_1 : boolean;
  signal call_stmt_846_call_ack_0 : boolean;
  signal slice_849_inst_ack_1 : boolean;
  signal call_stmt_846_call_req_0 : boolean;
  signal slice_849_inst_req_0 : boolean;
  signal call_stmt_846_call_req_1 : boolean;
  signal slice_849_inst_req_1 : boolean;
  signal slice_849_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryWord_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 169) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= word_addr_base;
  word_addr_base_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(136 downto 73) <= offset;
  offset_buffer <= in_buffer_data_out(136 downto 73);
  in_buffer_data_in(168 downto 137) <= wword;
  wword_buffer <= in_buffer_data_out(168 downto 137);
  in_buffer_data_in(tag_length + 168 downto 169) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 168 downto 169);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 1,6 => 7);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 7);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= tag_update_enable & rwbar_update_enable & word_addr_base_update_enable & offset_update_enable & wword_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryWord_CP_1007_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryWord_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rword_buffer;
  rword <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryWord_CP_1007_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rword_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rword_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rword_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rword_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryWord_CP_1007_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryWord_CP_1007_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryWord_CP_1007: Block -- control-path 
    signal accessMemoryWord_CP_1007_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    accessMemoryWord_CP_1007_elements(0) <= accessMemoryWord_CP_1007_start;
    accessMemoryWord_CP_1007_symbol <= accessMemoryWord_CP_1007_elements(22);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_846_to_assign_stmt_850/$entry
      -- 
    accessMemoryWord_CP_1007_elements(1) <= accessMemoryWord_CP_1007_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_846_to_assign_stmt_850/tag_update_enable_out
      -- CP-element group 2: 	 call_stmt_846_to_assign_stmt_850/tag_update_enable
      -- 
    accessMemoryWord_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWord_CP_1007_elements(10);
      gj_accessMemoryWord_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	10 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_846_to_assign_stmt_850/rwbar_update_enable_out
      -- CP-element group 3: 	 call_stmt_846_to_assign_stmt_850/rwbar_update_enable
      -- 
    accessMemoryWord_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWord_CP_1007_elements(10);
      gj_accessMemoryWord_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	10 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	18 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_846_to_assign_stmt_850/word_addr_base_update_enable_out
      -- CP-element group 4: 	 call_stmt_846_to_assign_stmt_850/word_addr_base_update_enable
      -- 
    accessMemoryWord_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWord_CP_1007_elements(10);
      gj_accessMemoryWord_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_846_to_assign_stmt_850/offset_update_enable_out
      -- CP-element group 5: 	 call_stmt_846_to_assign_stmt_850/offset_update_enable
      -- 
    accessMemoryWord_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWord_CP_1007_elements(10);
      gj_accessMemoryWord_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	10 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	20 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 call_stmt_846_to_assign_stmt_850/wword_update_enable
      -- CP-element group 6: 	 call_stmt_846_to_assign_stmt_850/wword_update_enable_out
      -- 
    accessMemoryWord_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWord_CP_1007_elements(10);
      gj_accessMemoryWord_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 call_stmt_846_to_assign_stmt_850/rword_update_enable
      -- CP-element group 7: 	 call_stmt_846_to_assign_stmt_850/rword_update_enable_in
      -- 
    accessMemoryWord_CP_1007_elements(7) <= accessMemoryWord_CP_1007_elements(21);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_sample_start_
      -- CP-element group 8: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/$entry
      -- CP-element group 8: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/crr
      -- 
    crr_1032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWord_CP_1007_elements(8), ack => call_stmt_846_call_req_0); -- 
    accessMemoryWord_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWord_CP_1007_elements(1) & accessMemoryWord_CP_1007_elements(10);
      gj_accessMemoryWord_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_update_start_
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/ccr
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/$entry
      -- 
    ccr_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWord_CP_1007_elements(9), ack => call_stmt_846_call_req_1); -- 
    accessMemoryWord_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "accessMemoryWord_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWord_CP_1007_elements(11) & accessMemoryWord_CP_1007_elements(14);
      gj_accessMemoryWord_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: 	5 
    -- CP-element group 10: 	6 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/cra
      -- CP-element group 10: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/$exit
      -- CP-element group 10: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_sample_completed_
      -- 
    cra_1033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_846_call_ack_0, ack => accessMemoryWord_CP_1007_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/cca
      -- CP-element group 11: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/$exit
      -- CP-element group 11: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_update_completed_
      -- 
    cca_1038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_846_call_ack_1, ack => accessMemoryWord_CP_1007_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_846_to_assign_stmt_850/slice_849_Sample/$entry
      -- CP-element group 12: 	 call_stmt_846_to_assign_stmt_850/slice_849_sample_start_
      -- CP-element group 12: 	 call_stmt_846_to_assign_stmt_850/slice_849_Sample/rr
      -- 
    rr_1046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWord_CP_1007_elements(12), ack => slice_849_inst_req_0); -- 
    accessMemoryWord_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "accessMemoryWord_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWord_CP_1007_elements(11) & accessMemoryWord_CP_1007_elements(14);
      gj_accessMemoryWord_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_846_to_assign_stmt_850/slice_849_update_start_
      -- CP-element group 13: 	 call_stmt_846_to_assign_stmt_850/slice_849_Update/cr
      -- CP-element group 13: 	 call_stmt_846_to_assign_stmt_850/slice_849_Update/$entry
      -- 
    cr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWord_CP_1007_elements(13), ack => slice_849_inst_req_1); -- 
    accessMemoryWord_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "accessMemoryWord_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWord_CP_1007_elements(7) & accessMemoryWord_CP_1007_elements(15);
      gj_accessMemoryWord_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWord_CP_1007_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_846_to_assign_stmt_850/slice_849_Sample/$exit
      -- CP-element group 14: 	 call_stmt_846_to_assign_stmt_850/slice_849_sample_completed_
      -- CP-element group 14: 	 call_stmt_846_to_assign_stmt_850/slice_849_Sample/ra
      -- 
    ra_1047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_849_inst_ack_0, ack => accessMemoryWord_CP_1007_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (4) 
      -- CP-element group 15: 	 call_stmt_846_to_assign_stmt_850/slice_849_update_completed_
      -- CP-element group 15: 	 call_stmt_846_to_assign_stmt_850/slice_849_Update/ca
      -- CP-element group 15: 	 call_stmt_846_to_assign_stmt_850/slice_849_Update/$exit
      -- CP-element group 15: 	 call_stmt_846_to_assign_stmt_850/$exit
      -- 
    ca_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_849_inst_ack_1, ack => accessMemoryWord_CP_1007_elements(15)); -- 
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 tag_update_enable
      -- 
    accessMemoryWord_CP_1007_elements(16) <= accessMemoryWord_CP_1007_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rwbar_update_enable
      -- 
    accessMemoryWord_CP_1007_elements(17) <= accessMemoryWord_CP_1007_elements(3);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	4 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 word_addr_base_update_enable
      -- 
    accessMemoryWord_CP_1007_elements(18) <= accessMemoryWord_CP_1007_elements(4);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 offset_update_enable
      -- 
    accessMemoryWord_CP_1007_elements(19) <= accessMemoryWord_CP_1007_elements(5);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 wword_update_enable
      -- 
    accessMemoryWord_CP_1007_elements(20) <= accessMemoryWord_CP_1007_elements(6);
    -- CP-element group 21:  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	7 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 rword_update_enable
      -- 
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 $exit
      -- 
    accessMemoryWord_CP_1007_elements(22) <= accessMemoryWord_CP_1007_elements(15);
    --  hookup: inputs to control-path 
    accessMemoryWord_CP_1007_elements(21) <= rword_update_enable;
    -- hookup: output from control-path 
    wword_update_enable <= accessMemoryWord_CP_1007_elements(20);
    offset_update_enable <= accessMemoryWord_CP_1007_elements(19);
    word_addr_base_update_enable <= accessMemoryWord_CP_1007_elements(18);
    rwbar_update_enable <= accessMemoryWord_CP_1007_elements(17);
    tag_update_enable <= accessMemoryWord_CP_1007_elements(16);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u32_u64_844_wire : std_logic_vector(63 downto 0);
    signal MUX_838_wire : std_logic_vector(2 downto 0);
    signal R_LD_836_wire_constant : std_logic_vector(2 downto 0);
    signal R_ST_837_wire_constant : std_logic_vector(2 downto 0);
    signal rdword_846 : std_logic_vector(63 downto 0);
    signal type_cast_842_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_LD_836_wire_constant <= "100";
    R_ST_837_wire_constant <= "001";
    type_cast_842_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_838_inst
    MUX_838_wire <= R_LD_836_wire_constant when (rwbar_buffer(0) /=  '0') else R_ST_837_wire_constant;
    slice_849_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_849_inst_req_0;
      slice_849_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_849_inst_req_1;
      slice_849_inst_ack_1<= update_ack(0);
      slice_849_inst: SliceSplitProtocol generic map(name => "slice_849_inst", in_data_width => 64, high_index => 31, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdword_846, dout => rword_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow through binary operator CONCAT_u32_u64_844_inst
    process(type_cast_842_wire_constant, wword_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_842_wire_constant, wword_buffer, tmp_var);
      CONCAT_u32_u64_844_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_846_call 
    doMemAccess_call_group_0: Block -- 
      signal data_in: std_logic_vector(202 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 36);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_846_call_req_0;
      call_stmt_846_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_846_call_req_1;
      call_stmt_846_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      doMemAccess_call_group_0_gI: SplitGuardInterface generic map(name => "doMemAccess_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & MUX_838_wire & word_addr_base_buffer & offset_buffer & CONCAT_u32_u64_844_wire;
      rdword_846 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 203,
        owidth => 203,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => doMemAccess_call_reqs(0),
          ackR => doMemAccess_call_acks(0),
          dataR => doMemAccess_call_data(202 downto 0),
          tagR => doMemAccess_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => doMemAccess_return_acks(0), -- cross-over
          ackL => doMemAccess_return_reqs(0), -- cross-over
          dataL => doMemAccess_return_data(63 downto 0),
          tagL => doMemAccess_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemoryWord_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessMemoryWordBase is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    word_addr_base : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wword : in  std_logic_vector(31 downto 0);
    rword : out  std_logic_vector(31 downto 0);
    calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
    calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
    calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
    calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
    calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
    calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
    calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
    calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
    accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
    accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemoryWordBase;
architecture accessMemoryWordBase_arch of accessMemoryWordBase is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 170)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal word_addr_base_buffer :  std_logic_vector(63 downto 0);
  signal word_addr_base_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wword_buffer :  std_logic_vector(31 downto 0);
  signal wword_update_enable: Boolean;
  -- output port buffer signals
  signal rword_buffer :  std_logic_vector(31 downto 0);
  signal rword_update_enable: Boolean;
  signal accessMemoryWordBase_CP_506_start: Boolean;
  signal accessMemoryWordBase_CP_506_symbol: Boolean;
  -- volatile/operator module components. 
  component calculateAddress36 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      addr : out  std_logic_vector(35 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      request : in  std_logic_vector(109 downto 0);
      response : out  std_logic_vector(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_data : out  std_logic_vector(255 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_calculateAddress36_expr_503_inst_req_0 : boolean;
  signal call_calculateAddress36_expr_503_inst_ack_0 : boolean;
  signal call_calculateAddress36_expr_503_inst_req_1 : boolean;
  signal call_calculateAddress36_expr_503_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_521_inst_req_0 : boolean;
  signal CONCAT_u32_u64_521_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_521_inst_req_1 : boolean;
  signal CONCAT_u32_u64_521_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_527_inst_req_0 : boolean;
  signal CONCAT_u32_u64_527_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_527_inst_req_1 : boolean;
  signal CONCAT_u32_u64_527_inst_ack_1 : boolean;
  signal CONCAT_u1_u2_545_inst_req_0 : boolean;
  signal CONCAT_u1_u2_545_inst_ack_0 : boolean;
  signal CONCAT_u1_u2_545_inst_req_1 : boolean;
  signal CONCAT_u1_u2_545_inst_ack_1 : boolean;
  signal W_tag_518_delayed_3_0_556_inst_req_0 : boolean;
  signal W_tag_518_delayed_3_0_556_inst_ack_0 : boolean;
  signal W_tag_518_delayed_3_0_556_inst_req_1 : boolean;
  signal W_tag_518_delayed_3_0_556_inst_ack_1 : boolean;
  signal call_stmt_562_call_req_0 : boolean;
  signal call_stmt_562_call_ack_0 : boolean;
  signal call_stmt_562_call_req_1 : boolean;
  signal call_stmt_562_call_ack_1 : boolean;
  signal W_lw_535_delayed_11_0_571_inst_req_0 : boolean;
  signal W_lw_535_delayed_11_0_571_inst_ack_0 : boolean;
  signal W_lw_535_delayed_11_0_571_inst_req_1 : boolean;
  signal W_lw_535_delayed_11_0_571_inst_ack_1 : boolean;
  signal MUX_578_inst_req_0 : boolean;
  signal MUX_578_inst_ack_0 : boolean;
  signal MUX_578_inst_req_1 : boolean;
  signal MUX_578_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemoryWordBase_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 170) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= lock;
  lock_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(9 downto 9) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(9 downto 9);
  in_buffer_data_in(73 downto 10) <= word_addr_base;
  word_addr_base_buffer <= in_buffer_data_out(73 downto 10);
  in_buffer_data_in(137 downto 74) <= offset;
  offset_buffer <= in_buffer_data_out(137 downto 74);
  in_buffer_data_in(169 downto 138) <= wword;
  wword_buffer <= in_buffer_data_out(169 downto 138);
  in_buffer_data_in(tag_length + 169 downto 170) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 169 downto 170);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 1,7 => 7);
    constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1,7 => 7);
    constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 8); -- 
  begin -- 
    preds <= tag_update_enable & lock_update_enable & rwbar_update_enable & word_addr_base_update_enable & offset_update_enable & wword_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemoryWordBase_CP_506_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemoryWordBase_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rword_buffer;
  rword <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryWordBase_CP_506_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rword_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rword_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rword_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rword_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemoryWordBase_CP_506_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemoryWordBase_CP_506_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemoryWordBase_CP_506: Block -- control-path 
    signal accessMemoryWordBase_CP_506_elements: BooleanArray(48 downto 0);
    -- 
  begin -- 
    accessMemoryWordBase_CP_506_elements(0) <= accessMemoryWordBase_CP_506_start;
    accessMemoryWordBase_CP_506_symbol <= accessMemoryWordBase_CP_506_elements(48);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	21 
    -- CP-element group 1: 	25 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_504_to_assign_stmt_579/$entry
      -- 
    accessMemoryWordBase_CP_506_elements(1) <= accessMemoryWordBase_CP_506_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	27 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	41 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_504_to_assign_stmt_579/tag_update_enable
      -- CP-element group 2: 	 assign_stmt_504_to_assign_stmt_579/tag_update_enable_out
      -- 
    accessMemoryWordBase_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWordBase_CP_506_elements(27);
      gj_accessMemoryWordBase_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	23 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	42 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_504_to_assign_stmt_579/lock_update_enable_out
      -- CP-element group 3: 	 assign_stmt_504_to_assign_stmt_579/lock_update_enable
      -- 
    accessMemoryWordBase_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWordBase_CP_506_elements(23);
      gj_accessMemoryWordBase_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	23 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	43 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_504_to_assign_stmt_579/rwbar_update_enable
      -- CP-element group 4: 	 assign_stmt_504_to_assign_stmt_579/rwbar_update_enable_out
      -- 
    accessMemoryWordBase_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWordBase_CP_506_elements(23);
      gj_accessMemoryWordBase_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	44 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_504_to_assign_stmt_579/word_addr_base_update_enable
      -- CP-element group 5: 	 assign_stmt_504_to_assign_stmt_579/word_addr_base_update_enable_out
      -- 
    accessMemoryWordBase_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWordBase_CP_506_elements(11);
      gj_accessMemoryWordBase_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	45 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_504_to_assign_stmt_579/offset_update_enable
      -- CP-element group 6: 	 assign_stmt_504_to_assign_stmt_579/offset_update_enable_out
      -- 
    accessMemoryWordBase_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemoryWordBase_CP_506_elements(11);
      gj_accessMemoryWordBase_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	15 
    -- CP-element group 7: 	19 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	46 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_504_to_assign_stmt_579/wword_update_enable
      -- CP-element group 7: 	 assign_stmt_504_to_assign_stmt_579/wword_update_enable_out
      -- 
    accessMemoryWordBase_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(15) & accessMemoryWordBase_CP_506_elements(19);
      gj_accessMemoryWordBase_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	47 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	38 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 assign_stmt_504_to_assign_stmt_579/rword_update_enable_in
      -- CP-element group 8: 	 assign_stmt_504_to_assign_stmt_579/rword_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(8) <= accessMemoryWordBase_CP_506_elements(47);
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Sample/req
      -- CP-element group 9: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_sample_start_
      -- 
    req_533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(9), ack => call_calculateAddress36_expr_503_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "accessMemoryWordBase_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(1) & accessMemoryWordBase_CP_506_elements(11);
      gj_accessMemoryWordBase_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	31 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Update/$entry
      -- CP-element group 10: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_update_start_
      -- CP-element group 10: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Update/req
      -- 
    req_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(10), ack => call_calculateAddress36_expr_503_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(31) & accessMemoryWordBase_CP_506_elements(35) & accessMemoryWordBase_CP_506_elements(12);
      gj_accessMemoryWordBase_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Sample/ack
      -- CP-element group 11: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_sample_completed_
      -- 
    ack_534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_calculateAddress36_expr_503_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12: 	33 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_update_completed_
      -- CP-element group 12: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Update/$exit
      -- CP-element group 12: 	 assign_stmt_504_to_assign_stmt_579/call_calculateAddress36_expr_503_Update/ack
      -- 
    ack_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_calculateAddress36_expr_503_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_sample_start_
      -- CP-element group 13: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Sample/rr
      -- 
    rr_547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(13), ack => CONCAT_u32_u64_521_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(1) & accessMemoryWordBase_CP_506_elements(15);
      gj_accessMemoryWordBase_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	31 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_update_start_
      -- CP-element group 14: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Update/$entry
      -- CP-element group 14: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Update/cr
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(14), ack => CONCAT_u32_u64_521_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(16) & accessMemoryWordBase_CP_506_elements(31);
      gj_accessMemoryWordBase_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	7 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_sample_completed_
      -- CP-element group 15: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Sample/ra
      -- 
    ra_548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_521_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_update_completed_
      -- CP-element group 16: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Update/$exit
      -- CP-element group 16: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_521_Update/ca
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_521_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_sample_start_
      -- CP-element group 17: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Sample/rr
      -- 
    rr_561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(17), ack => CONCAT_u32_u64_527_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(1) & accessMemoryWordBase_CP_506_elements(19);
      gj_accessMemoryWordBase_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	31 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_update_start_
      -- CP-element group 18: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Update/$entry
      -- CP-element group 18: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Update/cr
      -- 
    cr_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(18), ack => CONCAT_u32_u64_527_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(20) & accessMemoryWordBase_CP_506_elements(31);
      gj_accessMemoryWordBase_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: 	7 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_sample_completed_
      -- CP-element group 19: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Sample/ra
      -- 
    ra_562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_527_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_update_completed_
      -- CP-element group 20: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Update/$exit
      -- CP-element group 20: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u32_u64_527_Update/ca
      -- 
    ca_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_527_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	1 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_sample_start_
      -- CP-element group 21: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Sample/rr
      -- 
    rr_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(21), ack => CONCAT_u1_u2_545_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(1) & accessMemoryWordBase_CP_506_elements(23);
      gj_accessMemoryWordBase_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: 	31 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_update_start_
      -- CP-element group 22: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Update/$entry
      -- CP-element group 22: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Update/cr
      -- 
    cr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(22), ack => CONCAT_u1_u2_545_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(24) & accessMemoryWordBase_CP_506_elements(31);
      gj_accessMemoryWordBase_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: 	3 
    -- CP-element group 23: 	4 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_sample_completed_
      -- CP-element group 23: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Sample/$exit
      -- CP-element group 23: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Sample/ra
      -- 
    ra_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u2_545_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_update_completed_
      -- CP-element group 24: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Update/$exit
      -- CP-element group 24: 	 assign_stmt_504_to_assign_stmt_579/CONCAT_u1_u2_545_Update/ca
      -- 
    ca_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u2_545_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	1 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_sample_start_
      -- CP-element group 25: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Sample/req
      -- 
    req_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(25), ack => W_tag_518_delayed_3_0_556_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(1) & accessMemoryWordBase_CP_506_elements(27);
      gj_accessMemoryWordBase_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: 	31 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_update_start_
      -- CP-element group 26: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Update/$entry
      -- CP-element group 26: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Update/req
      -- 
    req_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(26), ack => W_tag_518_delayed_3_0_556_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(28) & accessMemoryWordBase_CP_506_elements(31);
      gj_accessMemoryWordBase_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	2 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_sample_completed_
      -- CP-element group 27: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Sample/ack
      -- 
    ack_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_518_delayed_3_0_556_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_update_completed_
      -- CP-element group 28: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Update/$exit
      -- CP-element group 28: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_558_Update/ack
      -- 
    ack_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_518_delayed_3_0_556_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	12 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_sample_start_
      -- CP-element group 29: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Sample/$entry
      -- CP-element group 29: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Sample/crr
      -- 
    crr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(29), ack => call_stmt_562_call_req_0); -- 
    accessMemoryWordBase_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(16) & accessMemoryWordBase_CP_506_elements(20) & accessMemoryWordBase_CP_506_elements(24) & accessMemoryWordBase_CP_506_elements(28) & accessMemoryWordBase_CP_506_elements(12) & accessMemoryWordBase_CP_506_elements(31);
      gj_accessMemoryWordBase_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	39 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_update_start_
      -- CP-element group 30: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Update/$entry
      -- CP-element group 30: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Update/ccr
      -- 
    ccr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(30), ack => call_stmt_562_call_req_1); -- 
    accessMemoryWordBase_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(32) & accessMemoryWordBase_CP_506_elements(39);
      gj_accessMemoryWordBase_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	29 
    -- CP-element group 31: 	10 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_sample_completed_
      -- CP-element group 31: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Sample/cra
      -- 
    cra_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_562_call_ack_0, ack => accessMemoryWordBase_CP_506_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	37 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_update_completed_
      -- CP-element group 32: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Update/$exit
      -- CP-element group 32: 	 assign_stmt_504_to_assign_stmt_579/call_stmt_562_Update/cca
      -- 
    cca_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_562_call_ack_1, ack => accessMemoryWordBase_CP_506_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	12 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_sample_start_
      -- CP-element group 33: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Sample/$entry
      -- CP-element group 33: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Sample/req
      -- 
    req_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(33), ack => W_lw_535_delayed_11_0_571_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(12) & accessMemoryWordBase_CP_506_elements(35);
      gj_accessMemoryWordBase_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	39 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_update_start_
      -- CP-element group 34: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Update/$entry
      -- CP-element group 34: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Update/req
      -- 
    req_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(34), ack => W_lw_535_delayed_11_0_571_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(36) & accessMemoryWordBase_CP_506_elements(39);
      gj_accessMemoryWordBase_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_sample_completed_
      -- CP-element group 35: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Sample/ack
      -- 
    ack_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lw_535_delayed_11_0_571_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_update_completed_
      -- CP-element group 36: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Update/$exit
      -- CP-element group 36: 	 assign_stmt_504_to_assign_stmt_579/assign_stmt_573_Update/ack
      -- 
    ack_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lw_535_delayed_11_0_571_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	32 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_sample_start_
      -- CP-element group 37: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_start/$entry
      -- CP-element group 37: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_start/req
      -- 
    req_631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(37), ack => MUX_578_inst_req_0); -- 
    accessMemoryWordBase_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(32) & accessMemoryWordBase_CP_506_elements(36) & accessMemoryWordBase_CP_506_elements(39);
      gj_accessMemoryWordBase_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	8 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_update_start_
      -- CP-element group 38: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_complete/$entry
      -- CP-element group 38: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_complete/req
      -- 
    req_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemoryWordBase_CP_506_elements(38), ack => MUX_578_inst_req_1); -- 
    accessMemoryWordBase_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "accessMemoryWordBase_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemoryWordBase_CP_506_elements(8) & accessMemoryWordBase_CP_506_elements(40);
      gj_accessMemoryWordBase_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemoryWordBase_CP_506_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	30 
    -- CP-element group 39: 	34 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_sample_completed_
      -- CP-element group 39: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_start/$exit
      -- CP-element group 39: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_start/ack
      -- 
    ack_632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_578_inst_ack_0, ack => accessMemoryWordBase_CP_506_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	48 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 assign_stmt_504_to_assign_stmt_579/$exit
      -- CP-element group 40: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_update_completed_
      -- CP-element group 40: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_complete/$exit
      -- CP-element group 40: 	 assign_stmt_504_to_assign_stmt_579/MUX_578_complete/ack
      -- 
    ack_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_578_inst_ack_1, ack => accessMemoryWordBase_CP_506_elements(40)); -- 
    -- CP-element group 41:  place  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	2 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 tag_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(41) <= accessMemoryWordBase_CP_506_elements(2);
    -- CP-element group 42:  place  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	3 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 lock_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(42) <= accessMemoryWordBase_CP_506_elements(3);
    -- CP-element group 43:  place  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	4 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 rwbar_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(43) <= accessMemoryWordBase_CP_506_elements(4);
    -- CP-element group 44:  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	5 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 word_addr_base_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(44) <= accessMemoryWordBase_CP_506_elements(5);
    -- CP-element group 45:  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	6 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 offset_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(45) <= accessMemoryWordBase_CP_506_elements(6);
    -- CP-element group 46:  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	7 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 wword_update_enable
      -- 
    accessMemoryWordBase_CP_506_elements(46) <= accessMemoryWordBase_CP_506_elements(7);
    -- CP-element group 47:  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	8 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 rword_update_enable
      -- 
    -- CP-element group 48:  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	40 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 $exit
      -- 
    accessMemoryWordBase_CP_506_elements(48) <= accessMemoryWordBase_CP_506_elements(40);
    --  hookup: inputs to control-path 
    accessMemoryWordBase_CP_506_elements(47) <= rword_update_enable;
    -- hookup: output from control-path 
    tag_update_enable <= accessMemoryWordBase_CP_506_elements(41);
    lock_update_enable <= accessMemoryWordBase_CP_506_elements(42);
    rwbar_update_enable <= accessMemoryWordBase_CP_506_elements(43);
    word_addr_base_update_enable <= accessMemoryWordBase_CP_506_elements(44);
    offset_update_enable <= accessMemoryWordBase_CP_506_elements(45);
    wword_update_enable <= accessMemoryWordBase_CP_506_elements(46);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_510_510_delayed_3_0_546 : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_550_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u32_u64_493_493_delayed_3_0_522 : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_497_497_delayed_3_0_528 : std_logic_vector(63 downto 0);
    signal CONCAT_u36_u100_553_wire : std_logic_vector(99 downto 0);
    signal addr_dw_541 : std_logic_vector(35 downto 0);
    signal bmask_516 : std_logic_vector(7 downto 0);
    signal konst_507_wire_constant : std_logic_vector(35 downto 0);
    signal konst_514_wire_constant : std_logic_vector(7 downto 0);
    signal lw_509 : std_logic_vector(0 downto 0);
    signal lw_535_delayed_11_0_573 : std_logic_vector(0 downto 0);
    signal request_555 : std_logic_vector(109 downto 0);
    signal response_562 : std_logic_vector(64 downto 0);
    signal rhw_566 : std_logic_vector(31 downto 0);
    signal rlw_570 : std_logic_vector(31 downto 0);
    signal slice_537_wire : std_logic_vector(32 downto 0);
    signal tag_518_delayed_3_0_558 : std_logic_vector(7 downto 0);
    signal type_cast_513_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_526_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_539_wire_constant : std_logic_vector(2 downto 0);
    signal wdata_534 : std_logic_vector(63 downto 0);
    signal word_addr_504 : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    konst_507_wire_constant <= "000000000000000000000000000000000010";
    konst_514_wire_constant <= "11110000";
    type_cast_513_wire_constant <= "00001111";
    type_cast_519_wire_constant <= "00000000000000000000000000000000";
    type_cast_526_wire_constant <= "00000000000000000000000000000000";
    type_cast_539_wire_constant <= "000";
    -- flow-through select operator MUX_515_inst
    bmask_516 <= type_cast_513_wire_constant when (lw_509(0) /=  '0') else konst_514_wire_constant;
    -- flow-through select operator MUX_533_inst
    wdata_534 <= CONCAT_u32_u64_493_493_delayed_3_0_522 when (lw_509(0) /=  '0') else CONCAT_u32_u64_497_497_delayed_3_0_528;
    MUX_578_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_578_inst_req_0;
      MUX_578_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_578_inst_req_1;
      MUX_578_inst_ack_1<= update_ack(0);
      MUX_578_inst: SelectSplitProtocol generic map(name => "MUX_578_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => rlw_570, y => rhw_566, sel => lw_535_delayed_11_0_573, z => rword_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_537_inst
    slice_537_wire <= word_addr_504(35 downto 3);
    -- flow-through slice operator slice_565_inst
    rhw_566 <= response_562(63 downto 32);
    -- flow-through slice operator slice_569_inst
    rlw_570 <= response_562(31 downto 0);
    W_lw_535_delayed_11_0_571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lw_535_delayed_11_0_571_inst_req_0;
      W_lw_535_delayed_11_0_571_inst_ack_0<= wack(0);
      rreq(0) <= W_lw_535_delayed_11_0_571_inst_req_1;
      W_lw_535_delayed_11_0_571_inst_ack_1<= rack(0);
      W_lw_535_delayed_11_0_571_inst : InterlockBuffer generic map ( -- 
        name => "W_lw_535_delayed_11_0_571_inst",
        buffer_size => 11,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lw_509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lw_535_delayed_11_0_573,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_tag_518_delayed_3_0_556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_tag_518_delayed_3_0_556_inst_req_0;
      W_tag_518_delayed_3_0_556_inst_ack_0<= wack(0);
      rreq(0) <= W_tag_518_delayed_3_0_556_inst_req_1;
      W_tag_518_delayed_3_0_556_inst_ack_1<= rack(0);
      W_tag_518_delayed_3_0_556_inst : InterlockBuffer generic map ( -- 
        name => "W_tag_518_delayed_3_0_556_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_518_delayed_3_0_558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- flow through binary operator BITSEL_u36_u1_508_inst
    process(word_addr_504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(word_addr_504, konst_507_wire_constant, tmp_var);
      lw_509 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u10_u110_554_inst
    process(CONCAT_u2_u10_550_wire, CONCAT_u36_u100_553_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_550_wire, CONCAT_u36_u100_553_wire, tmp_var);
      request_555 <= tmp_var; --
    end process;
    -- shared split operator group (2) : CONCAT_u1_u2_545_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= lock_buffer & rwbar_buffer;
      CONCAT_u1_u2_510_510_delayed_3_0_546 <= data_out(1 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u2_545_inst_req_0;
      CONCAT_u1_u2_545_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u2_545_inst_req_1;
      CONCAT_u1_u2_545_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 2,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 3,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- flow through binary operator CONCAT_u2_u10_550_inst
    process(CONCAT_u1_u2_510_510_delayed_3_0_546, bmask_516) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_510_510_delayed_3_0_546, bmask_516, tmp_var);
      CONCAT_u2_u10_550_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : CONCAT_u32_u64_521_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_519_wire_constant & wword_buffer;
      CONCAT_u32_u64_493_493_delayed_3_0_522 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_521_inst_req_0;
      CONCAT_u32_u64_521_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_521_inst_req_1;
      CONCAT_u32_u64_521_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 3,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : CONCAT_u32_u64_527_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= wword_buffer;
      CONCAT_u32_u64_497_497_delayed_3_0_528 <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_527_inst_req_0;
      CONCAT_u32_u64_527_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_527_inst_req_1;
      CONCAT_u32_u64_527_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          buffering  => 3,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- flow through binary operator CONCAT_u33_u36_540_inst
    process(slice_537_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_537_wire, type_cast_539_wire_constant, tmp_var);
      addr_dw_541 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u36_u100_553_inst
    process(addr_dw_541, wdata_534) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_dw_541, wdata_534, tmp_var);
      CONCAT_u36_u100_553_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_calculateAddress36_expr_503_inst 
    calculateAddress36_call_group_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_calculateAddress36_expr_503_inst_req_0;
      call_calculateAddress36_expr_503_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_calculateAddress36_expr_503_inst_req_1;
      call_calculateAddress36_expr_503_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      calculateAddress36_call_group_0_gI: SplitGuardInterface generic map(name => "calculateAddress36_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= word_addr_base_buffer & offset_buffer;
      word_addr_504 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => calculateAddress36_call_reqs(0),
          ackR => calculateAddress36_call_acks(0),
          dataR => calculateAddress36_call_data(127 downto 0),
          tagR => calculateAddress36_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => calculateAddress36_return_acks(0), -- cross-over
          ackL => calculateAddress36_return_reqs(0), -- cross-over
          dataL => calculateAddress36_return_data(35 downto 0),
          tagL => calculateAddress36_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_562_call 
    accessMemoryBase_call_group_1: Block -- 
      signal data_in: std_logic_vector(117 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 11);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_562_call_req_0;
      call_stmt_562_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_562_call_req_1;
      call_stmt_562_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryBase_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryBase_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_518_delayed_3_0_558 & request_555;
      response_562 <= data_out(64 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 118,
        owidth => 118,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryBase_call_reqs(0),
          ackR => accessMemoryBase_call_acks(0),
          dataR => accessMemoryBase_call_data(117 downto 0),
          tagR => accessMemoryBase_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 65,
          owidth => 65,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryBase_return_acks(0), -- cross-over
          ackL => accessMemoryBase_return_reqs(0), -- cross-over
          dataL => accessMemoryBase_return_data(64 downto 0),
          tagL => accessMemoryBase_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end accessMemoryWordBase_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    base_addr : in  std_logic_vector(63 downto 0);
    index : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
    accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
    accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessQueueElement;
architecture accessQueueElement_arch of accessQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 169)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal base_addr_buffer :  std_logic_vector(63 downto 0);
  signal base_addr_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(31 downto 0);
  signal index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessQueueElement_CP_1517_start: Boolean;
  signal accessQueueElement_CP_1517_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1114_call_req_0 : boolean;
  signal call_stmt_1114_call_ack_0 : boolean;
  signal call_stmt_1114_call_ack_1 : boolean;
  signal call_stmt_1114_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessQueueElement_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 169) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= base_addr;
  base_addr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(104 downto 73) <= index;
  index_buffer <= in_buffer_data_out(104 downto 73);
  in_buffer_data_in(168 downto 105) <= wdata;
  wdata_buffer <= in_buffer_data_out(168 downto 105);
  in_buffer_data_in(tag_length + 168 downto 169) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 168 downto 169);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessQueueElement_CP_1517_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessQueueElement_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueElement_CP_1517_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessQueueElement_CP_1517_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueElement_CP_1517_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessQueueElement_CP_1517: Block -- control-path 
    signal accessQueueElement_CP_1517_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    accessQueueElement_CP_1517_elements(0) <= accessQueueElement_CP_1517_start;
    accessQueueElement_CP_1517_symbol <= accessQueueElement_CP_1517_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_update_start_
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_sample_start_
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/$entry
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Update/ccr
      -- 
    crr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueElement_CP_1517_elements(0), ack => call_stmt_1114_call_req_0); -- 
    ccr_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueElement_CP_1517_elements(0), ack => call_stmt_1114_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Sample/cra
      -- 
    cra_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1114_call_ack_0, ack => accessQueueElement_CP_1517_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_update_completed_
      -- CP-element group 2: 	 assign_stmt_1107_to_call_stmt_1114/$exit
      -- CP-element group 2: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Update/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1107_to_call_stmt_1114/call_stmt_1114_Update/cca
      -- 
    cca_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1114_call_ack_1, ack => accessQueueElement_CP_1517_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u29_u61_1103_wire : std_logic_vector(60 downto 0);
    signal offset_1107 : std_logic_vector(63 downto 0);
    signal type_cast_1101_wire_constant : std_logic_vector(28 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    type_cast_1101_wire_constant <= "00000000000000000000000000000";
    type_cast_1105_wire_constant <= "000";
    -- flow through binary operator CONCAT_u29_u61_1103_inst
    process(type_cast_1101_wire_constant, index_buffer) -- 
      variable tmp_var : std_logic_vector(60 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1101_wire_constant, index_buffer, tmp_var);
      CONCAT_u29_u61_1103_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u61_u64_1106_inst
    process(CONCAT_u29_u61_1103_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u29_u61_1103_wire, type_cast_1105_wire_constant, tmp_var);
      offset_1107 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1114_call 
    accessMemoryDword_call_group_0: Block -- 
      signal data_in: std_logic_vector(200 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1114_call_req_0;
      call_stmt_1114_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1114_call_req_1;
      call_stmt_1114_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDword_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rwbar_buffer & base_addr_buffer & offset_1107 & wdata_buffer;
      rdata_buffer <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 201,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(0),
          ackR => accessMemoryDword_call_acks(0),
          dataR => accessMemoryDword_call_data(200 downto 0),
          tagR => accessMemoryDword_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(0), -- cross-over
          ackL => accessMemoryDword_return_reqs(0), -- cross-over
          dataL => accessMemoryDword_return_data(63 downto 0),
          tagL => accessMemoryDword_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessQueueLength is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    qptr : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
    accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessQueueLength;
architecture accessQueueLength_arch of accessQueueLength is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 105)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessQueueLength_CP_1336_start: Boolean;
  signal accessQueueLength_CP_1336_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1000_call_req_0 : boolean;
  signal call_stmt_1000_call_ack_0 : boolean;
  signal call_stmt_1000_call_req_1 : boolean;
  signal call_stmt_1000_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessQueueLength_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 105) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= qptr;
  qptr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(104 downto 73) <= wdata;
  wdata_buffer <= in_buffer_data_out(104 downto 73);
  in_buffer_data_in(tag_length + 104 downto 105) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 104 downto 105);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessQueueLength_CP_1336_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessQueueLength_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueLength_CP_1336_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessQueueLength_CP_1336_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueLength_CP_1336_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessQueueLength_CP_1336: Block -- control-path 
    signal accessQueueLength_CP_1336_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    accessQueueLength_CP_1336_elements(0) <= accessQueueLength_CP_1336_start;
    accessQueueLength_CP_1336_symbol <= accessQueueLength_CP_1336_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1000/$entry
      -- CP-element group 0: 	 call_stmt_1000/call_stmt_1000_sample_start_
      -- CP-element group 0: 	 call_stmt_1000/call_stmt_1000_update_start_
      -- CP-element group 0: 	 call_stmt_1000/call_stmt_1000_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1000/call_stmt_1000_Sample/crr
      -- CP-element group 0: 	 call_stmt_1000/call_stmt_1000_Update/$entry
      -- CP-element group 0: 	 call_stmt_1000/call_stmt_1000_Update/ccr
      -- 
    crr_1349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueLength_CP_1336_elements(0), ack => call_stmt_1000_call_req_0); -- 
    ccr_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueLength_CP_1336_elements(0), ack => call_stmt_1000_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1000/call_stmt_1000_sample_completed_
      -- CP-element group 1: 	 call_stmt_1000/call_stmt_1000_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1000/call_stmt_1000_Sample/cra
      -- 
    cra_1350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1000_call_ack_0, ack => accessQueueLength_CP_1336_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1000/$exit
      -- CP-element group 2: 	 call_stmt_1000/call_stmt_1000_update_completed_
      -- CP-element group 2: 	 call_stmt_1000/call_stmt_1000_Update/$exit
      -- CP-element group 2: 	 call_stmt_1000/call_stmt_1000_Update/cca
      -- 
    cca_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1000_call_ack_1, ack => accessQueueLength_CP_1336_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_997_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_997_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001100";
    -- shared call operator group (0) : call_stmt_1000_call 
    accessMemoryWord_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1000_call_req_0;
      call_stmt_1000_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1000_call_req_1;
      call_stmt_1000_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWord_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryWord_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rwbar_buffer & qptr_buffer & konst_997_wire_constant & wdata_buffer;
      rdata_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWord_call_reqs(0),
          ackR => accessMemoryWord_call_acks(0),
          dataR => accessMemoryWord_call_data(168 downto 0),
          tagR => accessMemoryWord_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWord_return_acks(0), -- cross-over
          ackL => accessMemoryWord_return_reqs(0), -- cross-over
          dataL => accessMemoryWord_return_data(31 downto 0),
          tagL => accessMemoryWord_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessQueueLength_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessQueueMisc is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    qptr : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
    accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessQueueMisc;
architecture accessQueueMisc_arch of accessQueueMisc is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 105)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessQueueMisc_CP_1059_start: Boolean;
  signal accessQueueMisc_CP_1059_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_864_call_req_0 : boolean;
  signal call_stmt_864_call_ack_0 : boolean;
  signal call_stmt_864_call_req_1 : boolean;
  signal call_stmt_864_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessQueueMisc_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 105) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= qptr;
  qptr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(104 downto 73) <= wdata;
  wdata_buffer <= in_buffer_data_out(104 downto 73);
  in_buffer_data_in(tag_length + 104 downto 105) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 104 downto 105);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessQueueMisc_CP_1059_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessQueueMisc_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueMisc_CP_1059_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessQueueMisc_CP_1059_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueMisc_CP_1059_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessQueueMisc_CP_1059: Block -- control-path 
    signal accessQueueMisc_CP_1059_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    accessQueueMisc_CP_1059_elements(0) <= accessQueueMisc_CP_1059_start;
    accessQueueMisc_CP_1059_symbol <= accessQueueMisc_CP_1059_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_864/call_stmt_864_Sample/$entry
      -- CP-element group 0: 	 call_stmt_864/$entry
      -- CP-element group 0: 	 call_stmt_864/call_stmt_864_Sample/crr
      -- CP-element group 0: 	 call_stmt_864/call_stmt_864_update_start_
      -- CP-element group 0: 	 call_stmt_864/call_stmt_864_sample_start_
      -- CP-element group 0: 	 call_stmt_864/call_stmt_864_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_864/call_stmt_864_Update/ccr
      -- 
    crr_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueMisc_CP_1059_elements(0), ack => call_stmt_864_call_req_0); -- 
    ccr_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueMisc_CP_1059_elements(0), ack => call_stmt_864_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_864/call_stmt_864_Sample/$exit
      -- CP-element group 1: 	 call_stmt_864/call_stmt_864_sample_completed_
      -- CP-element group 1: 	 call_stmt_864/call_stmt_864_Sample/cra
      -- 
    cra_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_864_call_ack_0, ack => accessQueueMisc_CP_1059_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_864/call_stmt_864_Update/$exit
      -- CP-element group 2: 	 call_stmt_864/call_stmt_864_update_completed_
      -- CP-element group 2: 	 call_stmt_864/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_864/call_stmt_864_Update/cca
      -- 
    cca_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_864_call_ack_1, ack => accessQueueMisc_CP_1059_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_861_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_861_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011100";
    -- shared call operator group (0) : call_stmt_864_call 
    accessMemoryWord_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_864_call_req_0;
      call_stmt_864_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_864_call_req_1;
      call_stmt_864_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWord_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryWord_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rwbar_buffer & qptr_buffer & konst_861_wire_constant & wdata_buffer;
      rdata_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWord_call_reqs(0),
          ackR => accessMemoryWord_call_acks(0),
          dataR => accessMemoryWord_call_data(168 downto 0),
          tagR => accessMemoryWord_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWord_return_acks(0), -- cross-over
          ackL => accessMemoryWord_return_reqs(0), -- cross-over
          dataL => accessMemoryWord_return_data(31 downto 0),
          tagL => accessMemoryWord_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessQueueMisc_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessQueueReadIndex is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    qptr : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
    accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessQueueReadIndex;
architecture accessQueueReadIndex_arch of accessQueueReadIndex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 105)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessQueueReadIndex_CP_1262_start: Boolean;
  signal accessQueueReadIndex_CP_1262_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_952_call_req_0 : boolean;
  signal call_stmt_952_call_ack_0 : boolean;
  signal call_stmt_952_call_req_1 : boolean;
  signal call_stmt_952_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessQueueReadIndex_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 105) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= qptr;
  qptr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(104 downto 73) <= wdata;
  wdata_buffer <= in_buffer_data_out(104 downto 73);
  in_buffer_data_in(tag_length + 104 downto 105) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 104 downto 105);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessQueueReadIndex_CP_1262_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessQueueReadIndex_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueReadIndex_CP_1262_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessQueueReadIndex_CP_1262_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueReadIndex_CP_1262_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessQueueReadIndex_CP_1262: Block -- control-path 
    signal accessQueueReadIndex_CP_1262_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    accessQueueReadIndex_CP_1262_elements(0) <= accessQueueReadIndex_CP_1262_start;
    accessQueueReadIndex_CP_1262_symbol <= accessQueueReadIndex_CP_1262_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_952/$entry
      -- CP-element group 0: 	 call_stmt_952/call_stmt_952_sample_start_
      -- CP-element group 0: 	 call_stmt_952/call_stmt_952_update_start_
      -- CP-element group 0: 	 call_stmt_952/call_stmt_952_Sample/$entry
      -- CP-element group 0: 	 call_stmt_952/call_stmt_952_Sample/crr
      -- CP-element group 0: 	 call_stmt_952/call_stmt_952_Update/$entry
      -- CP-element group 0: 	 call_stmt_952/call_stmt_952_Update/ccr
      -- 
    crr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueReadIndex_CP_1262_elements(0), ack => call_stmt_952_call_req_0); -- 
    ccr_1280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueReadIndex_CP_1262_elements(0), ack => call_stmt_952_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_952/call_stmt_952_sample_completed_
      -- CP-element group 1: 	 call_stmt_952/call_stmt_952_Sample/$exit
      -- CP-element group 1: 	 call_stmt_952/call_stmt_952_Sample/cra
      -- 
    cra_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_952_call_ack_0, ack => accessQueueReadIndex_CP_1262_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_952/$exit
      -- CP-element group 2: 	 call_stmt_952/call_stmt_952_update_completed_
      -- CP-element group 2: 	 call_stmt_952/call_stmt_952_Update/$exit
      -- CP-element group 2: 	 call_stmt_952/call_stmt_952_Update/cca
      -- 
    cca_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_952_call_ack_1, ack => accessQueueReadIndex_CP_1262_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_949_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_949_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    -- shared call operator group (0) : call_stmt_952_call 
    accessMemoryWord_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_952_call_req_0;
      call_stmt_952_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_952_call_req_1;
      call_stmt_952_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWord_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryWord_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rwbar_buffer & qptr_buffer & konst_949_wire_constant & wdata_buffer;
      rdata_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWord_call_reqs(0),
          ackR => accessMemoryWord_call_acks(0),
          dataR => accessMemoryWord_call_data(168 downto 0),
          tagR => accessMemoryWord_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWord_return_acks(0), -- cross-over
          ackL => accessMemoryWord_return_reqs(0), -- cross-over
          dataL => accessMemoryWord_return_data(31 downto 0),
          tagL => accessMemoryWord_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessQueueReadIndex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessQueueTotalMsgs is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    qptr : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
    accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessQueueTotalMsgs;
architecture accessQueueTotalMsgs_arch of accessQueueTotalMsgs is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 105)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessQueueTotalMsgs_CP_1376_start: Boolean;
  signal accessQueueTotalMsgs_CP_1376_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1026_call_req_0 : boolean;
  signal call_stmt_1026_call_ack_0 : boolean;
  signal call_stmt_1026_call_req_1 : boolean;
  signal call_stmt_1026_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessQueueTotalMsgs_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 105) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= qptr;
  qptr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(104 downto 73) <= wdata;
  wdata_buffer <= in_buffer_data_out(104 downto 73);
  in_buffer_data_in(tag_length + 104 downto 105) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 104 downto 105);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessQueueTotalMsgs_CP_1376_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessQueueTotalMsgs_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueTotalMsgs_CP_1376_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessQueueTotalMsgs_CP_1376_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueTotalMsgs_CP_1376_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessQueueTotalMsgs_CP_1376: Block -- control-path 
    signal accessQueueTotalMsgs_CP_1376_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    accessQueueTotalMsgs_CP_1376_elements(0) <= accessQueueTotalMsgs_CP_1376_start;
    accessQueueTotalMsgs_CP_1376_symbol <= accessQueueTotalMsgs_CP_1376_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1026/$entry
      -- CP-element group 0: 	 call_stmt_1026/call_stmt_1026_sample_start_
      -- CP-element group 0: 	 call_stmt_1026/call_stmt_1026_update_start_
      -- CP-element group 0: 	 call_stmt_1026/call_stmt_1026_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1026/call_stmt_1026_Sample/crr
      -- CP-element group 0: 	 call_stmt_1026/call_stmt_1026_Update/$entry
      -- CP-element group 0: 	 call_stmt_1026/call_stmt_1026_Update/ccr
      -- 
    crr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueTotalMsgs_CP_1376_elements(0), ack => call_stmt_1026_call_req_0); -- 
    ccr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueTotalMsgs_CP_1376_elements(0), ack => call_stmt_1026_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1026/call_stmt_1026_sample_completed_
      -- CP-element group 1: 	 call_stmt_1026/call_stmt_1026_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1026/call_stmt_1026_Sample/cra
      -- 
    cra_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1026_call_ack_0, ack => accessQueueTotalMsgs_CP_1376_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1026/$exit
      -- CP-element group 2: 	 call_stmt_1026/call_stmt_1026_update_completed_
      -- CP-element group 2: 	 call_stmt_1026/call_stmt_1026_Update/$exit
      -- CP-element group 2: 	 call_stmt_1026/call_stmt_1026_Update/cca
      -- 
    cca_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1026_call_ack_1, ack => accessQueueTotalMsgs_CP_1376_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_1023_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1023_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_1026_call 
    accessMemoryWord_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1026_call_req_0;
      call_stmt_1026_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1026_call_req_1;
      call_stmt_1026_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWord_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryWord_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rwbar_buffer & qptr_buffer & konst_1023_wire_constant & wdata_buffer;
      rdata_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWord_call_reqs(0),
          ackR => accessMemoryWord_call_acks(0),
          dataR => accessMemoryWord_call_data(168 downto 0),
          tagR => accessMemoryWord_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWord_return_acks(0), -- cross-over
          ackL => accessMemoryWord_return_reqs(0), -- cross-over
          dataL => accessMemoryWord_return_data(31 downto 0),
          tagL => accessMemoryWord_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessQueueTotalMsgs_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessQueueWriteIndex is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    qptr : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
    accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessQueueWriteIndex;
architecture accessQueueWriteIndex_arch of accessQueueWriteIndex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 105)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessQueueWriteIndex_CP_1282_start: Boolean;
  signal accessQueueWriteIndex_CP_1282_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_966_call_req_0 : boolean;
  signal call_stmt_966_call_ack_0 : boolean;
  signal call_stmt_966_call_req_1 : boolean;
  signal call_stmt_966_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessQueueWriteIndex_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 105) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(8 downto 8) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(8 downto 8);
  in_buffer_data_in(72 downto 9) <= qptr;
  qptr_buffer <= in_buffer_data_out(72 downto 9);
  in_buffer_data_in(104 downto 73) <= wdata;
  wdata_buffer <= in_buffer_data_out(104 downto 73);
  in_buffer_data_in(tag_length + 104 downto 105) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 104 downto 105);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessQueueWriteIndex_CP_1282_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessQueueWriteIndex_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueWriteIndex_CP_1282_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessQueueWriteIndex_CP_1282_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessQueueWriteIndex_CP_1282_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessQueueWriteIndex_CP_1282: Block -- control-path 
    signal accessQueueWriteIndex_CP_1282_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    accessQueueWriteIndex_CP_1282_elements(0) <= accessQueueWriteIndex_CP_1282_start;
    accessQueueWriteIndex_CP_1282_symbol <= accessQueueWriteIndex_CP_1282_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_966/$entry
      -- CP-element group 0: 	 call_stmt_966/call_stmt_966_sample_start_
      -- CP-element group 0: 	 call_stmt_966/call_stmt_966_update_start_
      -- CP-element group 0: 	 call_stmt_966/call_stmt_966_Sample/$entry
      -- CP-element group 0: 	 call_stmt_966/call_stmt_966_Sample/crr
      -- CP-element group 0: 	 call_stmt_966/call_stmt_966_Update/$entry
      -- CP-element group 0: 	 call_stmt_966/call_stmt_966_Update/ccr
      -- 
    crr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueWriteIndex_CP_1282_elements(0), ack => call_stmt_966_call_req_0); -- 
    ccr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessQueueWriteIndex_CP_1282_elements(0), ack => call_stmt_966_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_966/call_stmt_966_sample_completed_
      -- CP-element group 1: 	 call_stmt_966/call_stmt_966_Sample/$exit
      -- CP-element group 1: 	 call_stmt_966/call_stmt_966_Sample/cra
      -- 
    cra_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_966_call_ack_0, ack => accessQueueWriteIndex_CP_1282_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_966/$exit
      -- CP-element group 2: 	 call_stmt_966/call_stmt_966_update_completed_
      -- CP-element group 2: 	 call_stmt_966/call_stmt_966_Update/$exit
      -- CP-element group 2: 	 call_stmt_966/call_stmt_966_Update/cca
      -- 
    cca_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_966_call_ack_1, ack => accessQueueWriteIndex_CP_1282_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_963_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_963_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    -- shared call operator group (0) : call_stmt_966_call 
    accessMemoryWord_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_966_call_req_0;
      call_stmt_966_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_966_call_req_1;
      call_stmt_966_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWord_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryWord_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rwbar_buffer & qptr_buffer & konst_963_wire_constant & wdata_buffer;
      rdata_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWord_call_reqs(0),
          ackR => accessMemoryWord_call_acks(0),
          dataR => accessMemoryWord_call_data(168 downto 0),
          tagR => accessMemoryWord_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWord_return_acks(0), -- cross-over
          ackL => accessMemoryWord_return_reqs(0), -- cross-over
          dataL => accessMemoryWord_return_data(31 downto 0),
          tagL => accessMemoryWord_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accessQueueWriteIndex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity accessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    index : in  std_logic_vector(7 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessRegister;
architecture accessRegister_arch of accessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 45)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessRegister_CP_3_start: Boolean;
  signal accessRegister_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_166_load_0_req_0 : boolean;
  signal array_obj_ref_166_load_0_ack_0 : boolean;
  signal array_obj_ref_166_load_0_req_1 : boolean;
  signal array_obj_ref_166_load_0_ack_1 : boolean;
  signal array_obj_ref_239_store_0_req_0 : boolean;
  signal array_obj_ref_239_store_0_ack_0 : boolean;
  signal array_obj_ref_239_store_0_req_1 : boolean;
  signal array_obj_ref_239_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 45) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(12 downto 5) <= index;
  index_buffer <= in_buffer_data_out(12 downto 5);
  in_buffer_data_in(44 downto 13) <= wdata;
  wdata_buffer <= in_buffer_data_out(44 downto 13);
  in_buffer_data_in(tag_length + 44 downto 45) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 44 downto 45);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessRegister_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessRegister_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessRegister_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessRegister_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessRegister_CP_3: Block -- control-path 
    signal accessRegister_CP_3_elements: BooleanArray(6 downto 0);
    -- 
  begin -- 
    accessRegister_CP_3_elements(0) <= accessRegister_CP_3_start;
    accessRegister_CP_3_symbol <= accessRegister_CP_3_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	5 
    -- CP-element group 0:  members (69) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_sample_start_
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_update_start_
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_offset_calculated
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_resized_0
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_computed_0
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_update_start_
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_offset_calculated
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_resized_0
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_computed_0
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/word_access_complete/word_0/cr
      -- 
    cr_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessRegister_CP_3_elements(0), ack => array_obj_ref_166_load_0_req_1); -- 
    rr_53_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_53_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessRegister_CP_3_elements(0), ack => array_obj_ref_166_load_0_req_0); -- 
    cr_131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessRegister_CP_3_elements(0), ack => array_obj_ref_239_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_sample_completed_
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Sample/word_access_start/word_0/ra
      -- 
    ra_54_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_166_load_0_ack_0, ack => accessRegister_CP_3_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_update_completed_
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/$exit
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/array_obj_ref_166_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/array_obj_ref_166_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/array_obj_ref_166_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_Update/array_obj_ref_166_Merge/merge_ack
      -- 
    ca_65_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_166_load_0_ack_1, ack => accessRegister_CP_3_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: 	6 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_sample_start_
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/array_obj_ref_239_Split/$entry
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/array_obj_ref_239_Split/$exit
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/array_obj_ref_239_Split/split_req
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/array_obj_ref_239_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/word_access_start/word_0/rr
      -- 
    rr_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessRegister_CP_3_elements(3), ack => array_obj_ref_239_store_0_req_0); -- 
    accessRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "accessRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessRegister_CP_3_elements(0) & accessRegister_CP_3_elements(2) & accessRegister_CP_3_elements(6);
      gj_accessRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessRegister_CP_3_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_sample_completed_
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Sample/word_access_start/word_0/ra
      -- 
    ra_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_239_store_0_ack_0, ack => accessRegister_CP_3_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_241/$exit
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_update_completed_
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/$exit
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_239_Update/word_access_complete/word_0/ca
      -- 
    ca_132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_239_store_0_ack_1, ack => accessRegister_CP_3_elements(5)); -- 
    -- CP-element group 6:  transition  delay-element  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	3 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 assign_stmt_167_to_assign_stmt_241/array_obj_ref_166_array_obj_ref_239_delay
      -- 
    -- Element group accessRegister_CP_3_elements(6) is a control-delay.
    cp_element_6_delay: control_delay_element  generic map(name => " 6_delay", delay_value => 1)  port map(req => accessRegister_CP_3_elements(1), ack => accessRegister_CP_3_elements(6), clk => clk, reset =>reset);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_225_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_234_wire : std_logic_vector(15 downto 0);
    signal MUX_220_wire : std_logic_vector(7 downto 0);
    signal MUX_224_wire : std_logic_vector(7 downto 0);
    signal MUX_229_wire : std_logic_vector(7 downto 0);
    signal MUX_233_wire : std_logic_vector(7 downto 0);
    signal R_index_165_resized : std_logic_vector(7 downto 0);
    signal R_index_165_scaled : std_logic_vector(7 downto 0);
    signal R_index_238_resized : std_logic_vector(7 downto 0);
    signal R_index_238_scaled : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_166_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_166_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_239_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_239_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_239_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_239_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_239_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_239_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_239_word_offset_0 : std_logic_vector(7 downto 0);
    signal b0_171 : std_logic_vector(0 downto 0);
    signal b1_175 : std_logic_vector(0 downto 0);
    signal b2_179 : std_logic_vector(0 downto 0);
    signal b3_183 : std_logic_vector(0 downto 0);
    signal r0_187 : std_logic_vector(7 downto 0);
    signal r1_191 : std_logic_vector(7 downto 0);
    signal r2_195 : std_logic_vector(7 downto 0);
    signal r3_199 : std_logic_vector(7 downto 0);
    signal w0_203 : std_logic_vector(7 downto 0);
    signal w1_207 : std_logic_vector(7 downto 0);
    signal w2_211 : std_logic_vector(7 downto 0);
    signal w3_215 : std_logic_vector(7 downto 0);
    signal wval_236 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_166_offset_scale_factor_0 <= "00000001";
    array_obj_ref_166_resized_base_address <= "00000000";
    array_obj_ref_166_word_offset_0 <= "00000000";
    array_obj_ref_239_offset_scale_factor_0 <= "00000001";
    array_obj_ref_239_resized_base_address <= "00000000";
    array_obj_ref_239_word_offset_0 <= "00000000";
    -- flow-through select operator MUX_220_inst
    MUX_220_wire <= w0_203 when (b0_171(0) /=  '0') else r0_187;
    -- flow-through select operator MUX_224_inst
    MUX_224_wire <= w1_207 when (b1_175(0) /=  '0') else r1_191;
    -- flow-through select operator MUX_229_inst
    MUX_229_wire <= w2_211 when (b2_179(0) /=  '0') else r2_195;
    -- flow-through select operator MUX_233_inst
    MUX_233_wire <= w3_215 when (b3_183(0) /=  '0') else r3_199;
    -- flow-through slice operator slice_170_inst
    b0_171 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_174_inst
    b1_175 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_178_inst
    b2_179 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_182_inst
    b3_183 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_186_inst
    r0_187 <= rdata_buffer(31 downto 24);
    -- flow-through slice operator slice_190_inst
    r1_191 <= rdata_buffer(23 downto 16);
    -- flow-through slice operator slice_194_inst
    r2_195 <= rdata_buffer(15 downto 8);
    -- flow-through slice operator slice_198_inst
    r3_199 <= rdata_buffer(7 downto 0);
    -- flow-through slice operator slice_202_inst
    w0_203 <= wdata_buffer(31 downto 24);
    -- flow-through slice operator slice_206_inst
    w1_207 <= wdata_buffer(23 downto 16);
    -- flow-through slice operator slice_210_inst
    w2_211 <= wdata_buffer(15 downto 8);
    -- flow-through slice operator slice_214_inst
    w3_215 <= wdata_buffer(7 downto 0);
    -- equivalence array_obj_ref_166_addr_0
    process(array_obj_ref_166_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_166_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_166_gather_scatter
    process(array_obj_ref_166_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_data_0;
      ov(31 downto 0) := iv;
      rdata_buffer <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_166_index_0_rename
    process(R_index_165_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_165_resized;
      ov(7 downto 0) := iv;
      R_index_165_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_166_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(7 downto 0) := iv;
      R_index_165_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_166_index_offset
    process(R_index_165_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_165_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_166_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_166_root_address_inst
    process(array_obj_ref_166_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_166_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_166_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_239_addr_0
    process(array_obj_ref_239_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_239_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_239_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_239_gather_scatter
    process(wval_236) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_236;
      ov(31 downto 0) := iv;
      array_obj_ref_239_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_239_index_0_rename
    process(R_index_238_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_238_resized;
      ov(7 downto 0) := iv;
      R_index_238_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_239_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(7 downto 0) := iv;
      R_index_238_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_239_index_offset
    process(R_index_238_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_238_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_239_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_239_root_address_inst
    process(array_obj_ref_239_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_239_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_239_root_address <= ov(7 downto 0);
      --
    end process;
    -- flow through binary operator CONCAT_u16_u32_235_inst
    process(CONCAT_u8_u16_225_wire, CONCAT_u8_u16_234_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_225_wire, CONCAT_u8_u16_234_wire, tmp_var);
      wval_236 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_225_inst
    process(MUX_220_wire, MUX_224_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_220_wire, MUX_224_wire, tmp_var);
      CONCAT_u8_u16_225_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_234_inst
    process(MUX_229_wire, MUX_233_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_229_wire, MUX_233_wire, tmp_var);
      CONCAT_u8_u16_234_wire <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_166_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_166_load_0_req_0;
      array_obj_ref_166_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_166_load_0_req_1;
      array_obj_ref_166_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_166_word_address_0;
      array_obj_ref_166_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(7 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : array_obj_ref_239_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_239_store_0_req_0;
      array_obj_ref_239_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_239_store_0_req_1;
      array_obj_ref_239_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_239_word_address_0;
      data_in <= array_obj_ref_239_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(7 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity acquireLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    lock_address_pointer : in  std_logic_vector(63 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemoryLdStub_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryLdStub_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryLdStub_call_data : out  std_logic_vector(135 downto 0);
    accessMemoryLdStub_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryLdStub_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryLdStub_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryLdStub_return_data : in   std_logic_vector(7 downto 0);
    accessMemoryLdStub_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireLock;
architecture acquireLock_arch of acquireLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal lock_address_pointer_buffer :  std_logic_vector(63 downto 0);
  signal lock_address_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireLock_CP_1176_start: Boolean;
  signal acquireLock_CP_1176_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryLdStub is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      byte_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      rbyte : out  std_logic_vector(7 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_927_call_ack_1 : boolean;
  signal call_stmt_927_call_ack_0 : boolean;
  signal if_stmt_928_branch_req_0 : boolean;
  signal call_stmt_927_call_req_1 : boolean;
  signal call_stmt_927_call_req_0 : boolean;
  signal if_stmt_928_branch_ack_1 : boolean;
  signal if_stmt_928_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= lock_address_pointer;
  lock_address_pointer_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireLock_CP_1176_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_1176_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireLock_CP_1176_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_1176_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireLock_CP_1176: Block -- control-path 
    signal acquireLock_CP_1176_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    acquireLock_CP_1176_elements(0) <= acquireLock_CP_1176_start;
    acquireLock_CP_1176_symbol <= acquireLock_CP_1176_elements(4);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_921/branch_block_stmt_921__entry__
      -- CP-element group 0: 	 branch_block_stmt_921/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/merge_stmt_922__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	5 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_sample_completed_
      -- 
    cra_1201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_927_call_ack_0, ack => acquireLock_CP_1176_elements(1)); -- 
    -- CP-element group 2:  branch  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	5 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Update/ca
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/EQ_u8_u1_931_inputs/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/EQ_u8_u1_931_inputs/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/EQ_u8_u1_931/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_eval_test/branch_req
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/EQ_u8_u1_931_place
      -- CP-element group 2: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_921/call_stmt_927/$exit
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928__entry__
      -- CP-element group 2: 	 branch_block_stmt_921/call_stmt_927__exit__
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_if_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/if_stmt_928_else_link/$entry
      -- 
    cca_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_927_call_ack_1, ack => acquireLock_CP_1176_elements(2)); -- 
    branch_req_1233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_1176_elements(2), ack => if_stmt_928_branch_req_0); -- 
    -- CP-element group 3:  transition  place  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	5 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_921/if_stmt_928_if_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_921/if_stmt_928_if_link/if_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_921/loopback
      -- CP-element group 3: 	 branch_block_stmt_921/loopback_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_921/loopback_PhiReq/$exit
      -- 
    if_choice_transition_1238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_928_branch_ack_1, ack => acquireLock_CP_1176_elements(3)); -- 
    -- CP-element group 4:  merge  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (8) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 branch_block_stmt_921/branch_block_stmt_921__exit__
      -- CP-element group 4: 	 branch_block_stmt_921/if_stmt_928__exit__
      -- CP-element group 4: 	 branch_block_stmt_921/$exit
      -- CP-element group 4: 	 branch_block_stmt_921/if_stmt_928_else_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_921/if_stmt_928_else_link/else_choice_transition
      -- CP-element group 4: 	 assign_stmt_938/$entry
      -- CP-element group 4: 	 assign_stmt_938/$exit
      -- 
    else_choice_transition_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_928_branch_ack_0, ack => acquireLock_CP_1176_elements(4)); -- 
    -- CP-element group 5:  merge  fork  transition  place  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: 	2 
    -- CP-element group 5:  members (13) 
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927__entry__
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Update/ccr
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Sample/crr
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_update_start_
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/call_stmt_927_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_921/call_stmt_927/$entry
      -- CP-element group 5: 	 branch_block_stmt_921/merge_stmt_922__exit__
      -- CP-element group 5: 	 branch_block_stmt_921/merge_stmt_922_PhiReqMerge
      -- CP-element group 5: 	 branch_block_stmt_921/merge_stmt_922_PhiAck/$entry
      -- CP-element group 5: 	 branch_block_stmt_921/merge_stmt_922_PhiAck/$exit
      -- CP-element group 5: 	 branch_block_stmt_921/merge_stmt_922_PhiAck/dummy
      -- 
    ccr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_1176_elements(5), ack => call_stmt_927_call_req_1); -- 
    crr_1200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_1176_elements(5), ack => call_stmt_927_call_req_0); -- 
    acquireLock_CP_1176_elements(5) <= OrReduce(acquireLock_CP_1176_elements(0) & acquireLock_CP_1176_elements(3));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_931_wire : std_logic_vector(0 downto 0);
    signal konst_925_wire_constant : std_logic_vector(63 downto 0);
    signal konst_930_wire_constant : std_logic_vector(7 downto 0);
    signal lock_val_927 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_925_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_930_wire_constant <= "11111111";
    if_stmt_928_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u8_u1_931_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_928_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_928_branch_req_0,
          ack0 => if_stmt_928_branch_ack_0,
          ack1 => if_stmt_928_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator EQ_u8_u1_931_inst
    process(lock_val_927) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(lock_val_927, konst_930_wire_constant, tmp_var);
      EQ_u8_u1_931_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_927_call 
    accessMemoryLdStub_call_group_0: Block -- 
      signal data_in: std_logic_vector(135 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_927_call_req_0;
      call_stmt_927_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_927_call_req_1;
      call_stmt_927_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryLdStub_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryLdStub_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & lock_address_pointer_buffer & konst_925_wire_constant;
      lock_val_927 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 136,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryLdStub_call_reqs(0),
          ackR => accessMemoryLdStub_call_acks(0),
          dataR => accessMemoryLdStub_call_data(135 downto 0),
          tagR => accessMemoryLdStub_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryLdStub_return_acks(0), -- cross-over
          ackL => accessMemoryLdStub_return_reqs(0), -- cross-over
          dataL => accessMemoryLdStub_return_data(7 downto 0),
          tagL => accessMemoryLdStub_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity calculateAddress36 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr_base : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    addr : out  std_logic_vector(35 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity calculateAddress36;
architecture calculateAddress36_arch of calculateAddress36 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_base_buffer :  std_logic_vector(63 downto 0);
  signal addr_base_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  -- output port buffer signals
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal calculateAddress36_CP_197_start: Boolean;
  signal calculateAddress36_CP_197_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ADD_u36_u36_283_inst_req_0 : boolean;
  signal ADD_u36_u36_283_inst_ack_0 : boolean;
  signal ADD_u36_u36_283_inst_req_1 : boolean;
  signal ADD_u36_u36_283_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "calculateAddress36_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr_base;
  addr_base_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= offset;
  offset_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 3) := (0 => 3,1 => 3,2 => 1,3 => 3);
    constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 3);
    constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 4); -- 
  begin -- 
    preds <= addr_base_update_enable & offset_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  calculateAddress36_CP_197_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "calculateAddress36_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= addr_buffer;
  addr <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 1,2 => 3);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= calculateAddress36_CP_197_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  addr_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "addr_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_addr_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => addr_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 3,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= calculateAddress36_CP_197_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= calculateAddress36_CP_197_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  calculateAddress36_CP_197: Block -- control-path 
    signal calculateAddress36_CP_197_elements: BooleanArray(12 downto 0);
    -- 
  begin -- 
    calculateAddress36_CP_197_elements(0) <= calculateAddress36_CP_197_start;
    calculateAddress36_CP_197_symbol <= calculateAddress36_CP_197_elements(12);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_284/$entry
      -- 
    calculateAddress36_CP_197_elements(1) <= calculateAddress36_CP_197_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_284/addr_base_update_enable
      -- CP-element group 2: 	 assign_stmt_284/addr_base_update_enable_out
      -- 
    calculateAddress36_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "calculateAddress36_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= calculateAddress36_CP_197_elements(7);
      gj_calculateAddress36_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => calculateAddress36_CP_197_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	7 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_284/offset_update_enable
      -- CP-element group 3: 	 assign_stmt_284/offset_update_enable_out
      -- 
    calculateAddress36_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "calculateAddress36_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= calculateAddress36_CP_197_elements(7);
      gj_calculateAddress36_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => calculateAddress36_CP_197_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	11 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_284/addr_update_enable
      -- CP-element group 4: 	 assign_stmt_284/addr_update_enable_in
      -- 
    calculateAddress36_CP_197_elements(4) <= calculateAddress36_CP_197_elements(11);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_284/ADD_u36_u36_283_sample_start_
      -- CP-element group 5: 	 assign_stmt_284/ADD_u36_u36_283_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_284/ADD_u36_u36_283_Sample/rr
      -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => calculateAddress36_CP_197_elements(5), ack => ADD_u36_u36_283_inst_req_0); -- 
    calculateAddress36_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "calculateAddress36_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= calculateAddress36_CP_197_elements(1) & calculateAddress36_CP_197_elements(7);
      gj_calculateAddress36_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => calculateAddress36_CP_197_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_284/ADD_u36_u36_283_update_start_
      -- CP-element group 6: 	 assign_stmt_284/ADD_u36_u36_283_Update/$entry
      -- CP-element group 6: 	 assign_stmt_284/ADD_u36_u36_283_Update/cr
      -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => calculateAddress36_CP_197_elements(6), ack => ADD_u36_u36_283_inst_req_1); -- 
    calculateAddress36_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "calculateAddress36_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= calculateAddress36_CP_197_elements(4) & calculateAddress36_CP_197_elements(8);
      gj_calculateAddress36_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => calculateAddress36_CP_197_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	3 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_284/ADD_u36_u36_283_sample_completed_
      -- CP-element group 7: 	 assign_stmt_284/ADD_u36_u36_283_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_284/ADD_u36_u36_283_Sample/ra
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_283_inst_ack_0, ack => calculateAddress36_CP_197_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (4) 
      -- CP-element group 8: 	 assign_stmt_284/$exit
      -- CP-element group 8: 	 assign_stmt_284/ADD_u36_u36_283_update_completed_
      -- CP-element group 8: 	 assign_stmt_284/ADD_u36_u36_283_Update/$exit
      -- CP-element group 8: 	 assign_stmt_284/ADD_u36_u36_283_Update/ca
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_283_inst_ack_1, ack => calculateAddress36_CP_197_elements(8)); -- 
    -- CP-element group 9:  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 addr_base_update_enable
      -- 
    calculateAddress36_CP_197_elements(9) <= calculateAddress36_CP_197_elements(2);
    -- CP-element group 10:  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 offset_update_enable
      -- 
    calculateAddress36_CP_197_elements(10) <= calculateAddress36_CP_197_elements(3);
    -- CP-element group 11:  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	4 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 addr_update_enable
      -- 
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 $exit
      -- 
    calculateAddress36_CP_197_elements(12) <= calculateAddress36_CP_197_elements(8);
    --  hookup: inputs to control-path 
    calculateAddress36_CP_197_elements(11) <= addr_update_enable;
    -- hookup: output from control-path 
    addr_base_update_enable <= calculateAddress36_CP_197_elements(9);
    offset_update_enable <= calculateAddress36_CP_197_elements(10);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal slice_280_wire : std_logic_vector(35 downto 0);
    signal slice_282_wire : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_280_inst
    slice_280_wire <= addr_base_buffer(35 downto 0);
    -- flow-through slice operator slice_282_inst
    slice_282_wire <= offset_buffer(35 downto 0);
    -- shared split operator group (0) : ADD_u36_u36_283_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_280_wire & slice_282_wire;
      addr_buffer <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_283_inst_req_0;
      ADD_u36_u36_283_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_283_inst_req_1;
      ADD_u36_u36_283_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 36, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- 
  end Block; -- data_path
  -- 
end calculateAddress36_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity controlDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    QUEUE_MONITOR_SIGNAL : in std_logic_vector(31 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    NIC_INTR_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_INTR_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_INTR_pipe_write_data : out  std_logic_vector(0 downto 0);
    NIC_INTR_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_INTR_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_INTR_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
    S_CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    S_CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    S_CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    S_NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    S_NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    S_NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    NIC_INTR_INTERNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_INTR_INTERNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_INTR_INTERNAL_pipe_write_data : out  std_logic_vector(0 downto 0);
    memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
    memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
    memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(1 downto 0);
    accessRegister_call_acks : in   std_logic_vector(1 downto 0);
    accessRegister_call_data : out  std_logic_vector(89 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(1 downto 0);
    accessRegister_return_acks : in   std_logic_vector(1 downto 0);
    accessRegister_return_data : in   std_logic_vector(63 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(3 downto 0);
    setGlobalSignals_call_reqs : out  std_logic_vector(0 downto 0);
    setGlobalSignals_call_acks : in   std_logic_vector(0 downto 0);
    setGlobalSignals_call_tag  :  out  std_logic_vector(0 downto 0);
    setGlobalSignals_return_reqs : out  std_logic_vector(0 downto 0);
    setGlobalSignals_return_acks : in   std_logic_vector(0 downto 0);
    setGlobalSignals_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity controlDaemon;
architecture controlDaemon_arch of controlDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal controlDaemon_CP_3762_start: Boolean;
  signal controlDaemon_CP_3762_symbol: Boolean;
  -- volatile/operator module components. 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setGlobalSignals is -- 
    generic (tag_length : integer); 
    port ( -- 
      NIC_INTR_ENABLE : in std_logic_vector(0 downto 0);
      NIC_INTR_INTERNAL : in std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_data : out  std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_memory_access_lock_2020_inst_req_1 : boolean;
  signal WPIPE_MAC_ENABLE_2029_inst_req_0 : boolean;
  signal WPIPE_NIC_INTR_2032_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2035_inst_req_0 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2035_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2035_inst_req_1 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2035_inst_ack_1 : boolean;
  signal WPIPE_NIC_INTR_2032_inst_req_1 : boolean;
  signal call_stmt_2028_call_req_1 : boolean;
  signal WPIPE_memory_access_lock_2020_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_2032_inst_req_0 : boolean;
  signal WPIPE_memory_access_lock_2020_inst_req_0 : boolean;
  signal call_stmt_2028_call_ack_0 : boolean;
  signal call_stmt_2028_call_ack_1 : boolean;
  signal WPIPE_MAC_ENABLE_2029_inst_ack_0 : boolean;
  signal call_stmt_2028_call_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_2029_inst_ack_1 : boolean;
  signal WPIPE_memory_access_lock_2020_inst_ack_1 : boolean;
  signal do_while_stmt_2049_branch_req_0 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_2041_inst_req_1 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_2041_inst_ack_1 : boolean;
  signal WPIPE_NIC_INTR_2032_inst_ack_1 : boolean;
  signal WPIPE_NIC_INTR_INTERNAL_2038_inst_ack_1 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_2044_inst_req_1 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_2044_inst_ack_1 : boolean;
  signal WPIPE_NIC_INTR_INTERNAL_2038_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_INTERNAL_2038_inst_req_1 : boolean;
  signal call_stmt_2091_call_req_1 : boolean;
  signal call_stmt_2091_call_ack_1 : boolean;
  signal WPIPE_NIC_INTR_INTERNAL_2038_inst_req_0 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_2041_inst_req_0 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_2041_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_2052_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_2052_inst_ack_0 : boolean;
  signal call_stmt_2091_call_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_2052_inst_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_2052_inst_ack_1 : boolean;
  signal call_stmt_2091_call_req_0 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_2044_inst_req_0 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_2044_inst_ack_0 : boolean;
  signal WPIPE_MAC_ENABLE_2029_inst_req_1 : boolean;
  signal call_stmt_2109_call_req_0 : boolean;
  signal call_stmt_2109_call_ack_0 : boolean;
  signal call_stmt_2109_call_req_1 : boolean;
  signal call_stmt_2109_call_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2116_inst_req_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2116_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2116_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2116_inst_ack_1 : boolean;
  signal do_while_stmt_2049_branch_ack_0 : boolean;
  signal do_while_stmt_2049_branch_ack_1 : boolean;
  signal W_ignq_2122_inst_req_0 : boolean;
  signal W_ignq_2122_inst_ack_0 : boolean;
  signal W_ignq_2122_inst_req_1 : boolean;
  signal W_ignq_2122_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "controlDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  controlDaemon_CP_3762_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "controlDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= controlDaemon_CP_3762_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= controlDaemon_CP_3762_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= controlDaemon_CP_3762_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  controlDaemon_CP_3762: Block -- control-path 
    signal controlDaemon_CP_3762_elements: BooleanArray(50 downto 0);
    -- 
  begin -- 
    controlDaemon_CP_3762_elements(0) <= controlDaemon_CP_3762_start;
    controlDaemon_CP_3762_symbol <= controlDaemon_CP_3762_elements(50);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_update_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Sample/req
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Sample/req
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Update/ccr
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Update/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Sample/req
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Sample/req
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Sample/crr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_sample_start_
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Sample/req
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Sample/req
      -- CP-element group 0: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Sample/req
      -- 
    req_3775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_memory_access_lock_2020_inst_req_0); -- 
    crr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => call_stmt_2028_call_req_0); -- 
    ccr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => call_stmt_2028_call_req_1); -- 
    req_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_MAC_ENABLE_2029_inst_req_0); -- 
    req_3817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_NIC_INTR_2032_inst_req_0); -- 
    req_3831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_NIC_INTR_ENABLE_2035_inst_req_0); -- 
    req_3845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_NIC_INTR_INTERNAL_2038_inst_req_0); -- 
    req_3859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_S_CONTROL_REGISTER_2041_inst_req_0); -- 
    req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(0), ack => WPIPE_S_NUMBER_OF_SERVERS_2044_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Update/req
      -- CP-element group 1: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_update_start_
      -- CP-element group 1: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Sample/ack
      -- CP-element group 1: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_sample_completed_
      -- CP-element group 1: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Update/$entry
      -- 
    ack_3776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_memory_access_lock_2020_inst_ack_0, ack => controlDaemon_CP_3762_elements(1)); -- 
    req_3780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(1), ack => WPIPE_memory_access_lock_2020_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_update_completed_
      -- CP-element group 2: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Update/$exit
      -- CP-element group 2: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_memory_access_lock_2020_Update/ack
      -- 
    ack_3781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_memory_access_lock_2020_inst_ack_1, ack => controlDaemon_CP_3762_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_sample_completed_
      -- CP-element group 3: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Sample/cra
      -- CP-element group 3: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Sample/$exit
      -- 
    cra_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2028_call_ack_0, ack => controlDaemon_CP_3762_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	17 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_update_completed_
      -- CP-element group 4: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Update/$exit
      -- CP-element group 4: 	 assign_stmt_2022_to_assign_stmt_2046/call_stmt_2028_Update/cca
      -- 
    cca_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2028_call_ack_1, ack => controlDaemon_CP_3762_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_update_start_
      -- CP-element group 5: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_sample_completed_
      -- CP-element group 5: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Update/$entry
      -- CP-element group 5: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Sample/ack
      -- CP-element group 5: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Update/req
      -- 
    ack_3804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_2029_inst_ack_0, ack => controlDaemon_CP_3762_elements(5)); -- 
    req_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(5), ack => WPIPE_MAC_ENABLE_2029_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	17 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_update_completed_
      -- CP-element group 6: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Update/$exit
      -- CP-element group 6: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_MAC_ENABLE_2029_Update/ack
      -- 
    ack_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_2029_inst_ack_1, ack => controlDaemon_CP_3762_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Update/$entry
      -- CP-element group 7: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Sample/ack
      -- CP-element group 7: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Update/req
      -- CP-element group 7: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_sample_completed_
      -- CP-element group 7: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_update_start_
      -- 
    ack_3818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_2032_inst_ack_0, ack => controlDaemon_CP_3762_elements(7)); -- 
    req_3822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(7), ack => WPIPE_NIC_INTR_2032_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	17 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Update/$exit
      -- CP-element group 8: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_Update/ack
      -- CP-element group 8: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_2032_update_completed_
      -- 
    ack_3823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_2032_inst_ack_1, ack => controlDaemon_CP_3762_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Update/$entry
      -- CP-element group 9: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Sample/ack
      -- CP-element group 9: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_update_start_
      -- CP-element group 9: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_sample_completed_
      -- CP-element group 9: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Update/req
      -- 
    ack_3832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_ENABLE_2035_inst_ack_0, ack => controlDaemon_CP_3762_elements(9)); -- 
    req_3836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(9), ack => WPIPE_NIC_INTR_ENABLE_2035_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	17 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Update/$exit
      -- CP-element group 10: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_update_completed_
      -- CP-element group 10: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_ENABLE_2035_Update/ack
      -- 
    ack_3837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_ENABLE_2035_inst_ack_1, ack => controlDaemon_CP_3762_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_update_start_
      -- CP-element group 11: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_sample_completed_
      -- CP-element group 11: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Sample/ack
      -- CP-element group 11: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Update/req
      -- CP-element group 11: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Update/$entry
      -- 
    ack_3846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_INTERNAL_2038_inst_ack_0, ack => controlDaemon_CP_3762_elements(11)); -- 
    req_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(11), ack => WPIPE_NIC_INTR_INTERNAL_2038_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	17 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_update_completed_
      -- CP-element group 12: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Update/ack
      -- CP-element group 12: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_NIC_INTR_INTERNAL_2038_Update/$exit
      -- 
    ack_3851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_INTERNAL_2038_inst_ack_1, ack => controlDaemon_CP_3762_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_sample_completed_
      -- CP-element group 13: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Update/req
      -- CP-element group 13: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_update_start_
      -- CP-element group 13: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Sample/ack
      -- CP-element group 13: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Update/$entry
      -- 
    ack_3860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_CONTROL_REGISTER_2041_inst_ack_0, ack => controlDaemon_CP_3762_elements(13)); -- 
    req_3864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(13), ack => WPIPE_S_CONTROL_REGISTER_2041_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Update/ack
      -- CP-element group 14: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_update_completed_
      -- CP-element group 14: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_CONTROL_REGISTER_2041_Update/$exit
      -- 
    ack_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_CONTROL_REGISTER_2041_inst_ack_1, ack => controlDaemon_CP_3762_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_update_start_
      -- CP-element group 15: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Update/$entry
      -- CP-element group 15: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Update/req
      -- CP-element group 15: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_sample_completed_
      -- CP-element group 15: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Sample/ack
      -- 
    ack_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_NUMBER_OF_SERVERS_2044_inst_ack_0, ack => controlDaemon_CP_3762_elements(15)); -- 
    req_3878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(15), ack => WPIPE_S_NUMBER_OF_SERVERS_2044_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_update_completed_
      -- CP-element group 16: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Update/$exit
      -- CP-element group 16: 	 assign_stmt_2022_to_assign_stmt_2046/WPIPE_S_NUMBER_OF_SERVERS_2044_Update/ack
      -- 
    ack_3879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_NUMBER_OF_SERVERS_2044_inst_ack_1, ack => controlDaemon_CP_3762_elements(16)); -- 
    -- CP-element group 17:  join  transition  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: 	4 
    -- CP-element group 17: 	6 
    -- CP-element group 17: 	8 
    -- CP-element group 17: 	10 
    -- CP-element group 17: 	12 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_2048/do_while_stmt_2049__entry__
      -- CP-element group 17: 	 branch_block_stmt_2048/$entry
      -- CP-element group 17: 	 assign_stmt_2022_to_assign_stmt_2046/$exit
      -- CP-element group 17: 	 branch_block_stmt_2048/branch_block_stmt_2048__entry__
      -- 
    controlDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(2) & controlDaemon_CP_3762_elements(4) & controlDaemon_CP_3762_elements(6) & controlDaemon_CP_3762_elements(8) & controlDaemon_CP_3762_elements(10) & controlDaemon_CP_3762_elements(12) & controlDaemon_CP_3762_elements(14) & controlDaemon_CP_3762_elements(16);
      gj_controlDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  place  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	48 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	49 
    -- CP-element group 18: 	50 
    -- CP-element group 18:  members (10) 
      -- CP-element group 18: 	 branch_block_stmt_2048/do_while_stmt_2049__exit__
      -- CP-element group 18: 	 branch_block_stmt_2048/$exit
      -- CP-element group 18: 	 branch_block_stmt_2048/branch_block_stmt_2048__exit__
      -- CP-element group 18: 	 assign_stmt_2124/$entry
      -- CP-element group 18: 	 assign_stmt_2124/assign_stmt_2124_sample_start_
      -- CP-element group 18: 	 assign_stmt_2124/assign_stmt_2124_update_start_
      -- CP-element group 18: 	 assign_stmt_2124/assign_stmt_2124_Sample/$entry
      -- CP-element group 18: 	 assign_stmt_2124/assign_stmt_2124_Sample/req
      -- CP-element group 18: 	 assign_stmt_2124/assign_stmt_2124_Update/$entry
      -- CP-element group 18: 	 assign_stmt_2124/assign_stmt_2124_Update/req
      -- 
    req_3982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(18), ack => W_ignq_2122_inst_req_0); -- 
    req_3987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(18), ack => W_ignq_2122_inst_req_1); -- 
    controlDaemon_CP_3762_elements(18) <= controlDaemon_CP_3762_elements(48);
    -- CP-element group 19:  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	25 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049__entry__
      -- CP-element group 19: 	 branch_block_stmt_2048/do_while_stmt_2049/$entry
      -- 
    controlDaemon_CP_3762_elements(19) <= controlDaemon_CP_3762_elements(17);
    -- CP-element group 20:  merge  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	48 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049__exit__
      -- 
    -- Element group controlDaemon_CP_3762_elements(20) is bound as output of CP function.
    -- CP-element group 21:  merge  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_back
      -- 
    -- Element group controlDaemon_CP_3762_elements(21) is bound as output of CP function.
    -- CP-element group 22:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	43 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	46 
    -- CP-element group 22: 	47 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2048/do_while_stmt_2049/condition_done
      -- CP-element group 22: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_exit/$entry
      -- CP-element group 22: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_taken/$entry
      -- 
    controlDaemon_CP_3762_elements(22) <= controlDaemon_CP_3762_elements(43);
    -- CP-element group 23:  branch  place  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	45 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_body_done
      -- 
    controlDaemon_CP_3762_elements(23) <= controlDaemon_CP_3762_elements(45);
    -- CP-element group 24:  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/back_edge_to_loop_body
      -- 
    controlDaemon_CP_3762_elements(24) <= controlDaemon_CP_3762_elements(21);
    -- CP-element group 25:  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	19 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/first_time_through_loop_body
      -- 
    controlDaemon_CP_3762_elements(25) <= controlDaemon_CP_3762_elements(19);
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	43 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/loop_body_start
      -- CP-element group 26: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/$entry
      -- 
    -- Element group controlDaemon_CP_3762_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Sample/rr
      -- 
    rr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(27), ack => RPIPE_AFB_NIC_REQUEST_2052_inst_req_0); -- 
    controlDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(26) & controlDaemon_CP_3762_elements(30);
      gj_controlDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	33 
    -- CP-element group 28: 	38 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Update/cr
      -- 
    cr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(28), ack => RPIPE_AFB_NIC_REQUEST_2052_inst_req_1); -- 
    controlDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(29) & controlDaemon_CP_3762_elements(33) & controlDaemon_CP_3762_elements(38);
      gj_controlDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Sample/ra
      -- 
    ra_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_2052_inst_ack_0, ack => controlDaemon_CP_3762_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	36 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/RPIPE_AFB_NIC_REQUEST_2052_Update/ca
      -- 
    ca_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_2052_inst_ack_1, ack => controlDaemon_CP_3762_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	39 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Sample/crr
      -- 
    crr_3924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(31), ack => call_stmt_2091_call_req_0); -- 
    controlDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(30) & controlDaemon_CP_3762_elements(33) & controlDaemon_CP_3762_elements(39);
      gj_controlDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: 	41 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Update/ccr
      -- CP-element group 32: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_update_start_
      -- 
    ccr_3929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(32), ack => call_stmt_2091_call_req_1); -- 
    controlDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(34) & controlDaemon_CP_3762_elements(41);
      gj_controlDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Sample/cra
      -- CP-element group 33: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Sample/$exit
      -- 
    cra_3925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2091_call_ack_0, ack => controlDaemon_CP_3762_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	44 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Update/cca
      -- CP-element group 34: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_update_completed_
      -- 
    cca_3930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2091_call_ack_1, ack => controlDaemon_CP_3762_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	40 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/barrier_stmt_2092_update_completed_
      -- 
    controlDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(30) & controlDaemon_CP_3762_elements(34);
      gj_controlDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	30 
    -- CP-element group 36: 	44 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Sample/crr
      -- 
    crr_3939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(36), ack => call_stmt_2109_call_req_0); -- 
    controlDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(30) & controlDaemon_CP_3762_elements(44) & controlDaemon_CP_3762_elements(38);
      gj_controlDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Update/ccr
      -- 
    ccr_3944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(37), ack => call_stmt_2109_call_req_1); -- 
    controlDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= controlDaemon_CP_3762_elements(39);
      gj_controlDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	28 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Sample/cra
      -- 
    cra_3940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2109_call_ack_0, ack => controlDaemon_CP_3762_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	45 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	31 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2109_Update/cca
      -- CP-element group 39: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/ring_reenable_memory_space_0
      -- 
    cca_3945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2109_call_ack_1, ack => controlDaemon_CP_3762_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: 	35 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Sample/req
      -- 
    req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(40), ack => WPIPE_AFB_NIC_RESPONSE_2116_inst_req_0); -- 
    controlDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(34) & controlDaemon_CP_3762_elements(35) & controlDaemon_CP_3762_elements(42);
      gj_controlDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	32 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_update_start_
      -- CP-element group 41: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Update/req
      -- 
    ack_3954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_2116_inst_ack_0, ack => controlDaemon_CP_3762_elements(41)); -- 
    req_3958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(41), ack => WPIPE_AFB_NIC_RESPONSE_2116_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/WPIPE_AFB_NIC_RESPONSE_2116_Update/ack
      -- 
    ack_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_2116_inst_ack_1, ack => controlDaemon_CP_3762_elements(42)); -- 
    -- CP-element group 43:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	26 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	22 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/condition_evaluated
      -- CP-element group 43: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_3901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => controlDaemon_CP_3762_elements(43), ack => do_while_stmt_2049_branch_req_0); -- 
    -- Element group controlDaemon_CP_3762_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => controlDaemon_CP_3762_elements(26), ack => controlDaemon_CP_3762_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	34 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	36 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/call_stmt_2091_call_stmt_2109_delay
      -- 
    -- Element group controlDaemon_CP_3762_elements(44) is a control-delay.
    cp_element_44_delay: control_delay_element  generic map(name => " 44_delay", delay_value => 1)  port map(req => controlDaemon_CP_3762_elements(34), ack => controlDaemon_CP_3762_elements(44), clk => clk, reset =>reset);
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	39 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	23 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_2048/do_while_stmt_2049/do_while_stmt_2049_loop_body/$exit
      -- 
    controlDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "controlDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= controlDaemon_CP_3762_elements(39) & controlDaemon_CP_3762_elements(42);
      gj_controlDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => controlDaemon_CP_3762_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	22 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_exit/$exit
      -- CP-element group 46: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_exit/ack
      -- 
    ack_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2049_branch_ack_0, ack => controlDaemon_CP_3762_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	22 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_taken/$exit
      -- CP-element group 47: 	 branch_block_stmt_2048/do_while_stmt_2049/loop_taken/ack
      -- 
    ack_3970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2049_branch_ack_1, ack => controlDaemon_CP_3762_elements(47)); -- 
    -- CP-element group 48:  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	20 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	18 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2048/do_while_stmt_2049/$exit
      -- 
    controlDaemon_CP_3762_elements(48) <= controlDaemon_CP_3762_elements(20);
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	18 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_2124/assign_stmt_2124_sample_completed_
      -- CP-element group 49: 	 assign_stmt_2124/assign_stmt_2124_Sample/$exit
      -- CP-element group 49: 	 assign_stmt_2124/assign_stmt_2124_Sample/ack
      -- 
    ack_3983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ignq_2122_inst_ack_0, ack => controlDaemon_CP_3762_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	18 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 $exit
      -- CP-element group 50: 	 assign_stmt_2124/$exit
      -- CP-element group 50: 	 assign_stmt_2124/assign_stmt_2124_update_completed_
      -- CP-element group 50: 	 assign_stmt_2124/assign_stmt_2124_Update/$exit
      -- CP-element group 50: 	 assign_stmt_2124/assign_stmt_2124_Update/ack
      -- 
    ack_3988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ignq_2122_inst_ack_1, ack => controlDaemon_CP_3762_elements(50)); -- 
    controlDaemon_do_while_stmt_2049_terminator_3971: loop_terminator -- 
      generic map (name => " controlDaemon_do_while_stmt_2049_terminator_3971", max_iterations_in_flight =>3) 
      port map(loop_body_exit => controlDaemon_CP_3762_elements(23),loop_continue => controlDaemon_CP_3762_elements(47),loop_terminate => controlDaemon_CP_3762_elements(46),loop_back => controlDaemon_CP_3762_elements(21),loop_exit => controlDaemon_CP_3762_elements(20),clk => clk, reset => reset); -- 
    entry_tmerge_3902_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= controlDaemon_CP_3762_elements(24);
        preds(1)  <= controlDaemon_CP_3762_elements(25);
        entry_tmerge_3902 : transition_merge -- 
          generic map(name => " entry_tmerge_3902")
          port map (preds => preds, symbol_out => controlDaemon_CP_3762_elements(26));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_2105_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_2098_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2095_wire : std_logic_vector(0 downto 0);
    signal RPIPE_QUEUE_MONITOR_SIGNAL_2123_wire : std_logic_vector(31 downto 0);
    signal addr_2071 : std_logic_vector(35 downto 0);
    signal bmask_2067 : std_logic_vector(3 downto 0);
    signal ign_2028 : std_logic_vector(31 downto 0);
    signal ignq_2124 : std_logic_vector(31 downto 0);
    signal index_2085 : std_logic_vector(7 downto 0);
    signal konst_2021_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2023_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2024_wire_constant : std_logic_vector(3 downto 0);
    signal konst_2025_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2026_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2030_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2033_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2036_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2039_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2042_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2045_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2097_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2104_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2120_wire_constant : std_logic_vector(0 downto 0);
    signal lock_2059 : std_logic_vector(0 downto 0);
    signal rdata_2091 : std_logic_vector(31 downto 0);
    signal req_2053 : std_logic_vector(73 downto 0);
    signal resp_2115 : std_logic_vector(32 downto 0);
    signal rwbar_2063 : std_logic_vector(0 downto 0);
    signal set_globals_2107 : std_logic_vector(0 downto 0);
    signal type_cast_2112_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_2100 : std_logic_vector(0 downto 0);
    signal wdata_2075 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_2021_wire_constant <= "1";
    konst_2023_wire_constant <= "0";
    konst_2024_wire_constant <= "0000";
    konst_2025_wire_constant <= "00000000";
    konst_2026_wire_constant <= "00000000000000000000000000000000";
    konst_2030_wire_constant <= "0";
    konst_2033_wire_constant <= "0";
    konst_2036_wire_constant <= "0";
    konst_2039_wire_constant <= "0";
    konst_2042_wire_constant <= "00000000000000000000000000000000";
    konst_2045_wire_constant <= "00000000000000000000000000000000";
    konst_2097_wire_constant <= "00000000";
    konst_2104_wire_constant <= "00000000000000000000000000000000";
    konst_2120_wire_constant <= "1";
    type_cast_2112_wire_constant <= "0";
    -- flow-through slice operator slice_2058_inst
    lock_2059 <= req_2053(73 downto 73);
    -- flow-through slice operator slice_2062_inst
    rwbar_2063 <= req_2053(72 downto 72);
    -- flow-through slice operator slice_2066_inst
    bmask_2067 <= req_2053(71 downto 68);
    -- flow-through slice operator slice_2070_inst
    addr_2071 <= req_2053(67 downto 32);
    -- flow-through slice operator slice_2074_inst
    wdata_2075 <= req_2053(31 downto 0);
    -- flow-through slice operator slice_2084_inst
    index_2085 <= addr_2071(9 downto 2);
    W_ignq_2122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ignq_2122_inst_req_0;
      W_ignq_2122_inst_ack_0<= wack(0);
      rreq(0) <= W_ignq_2122_inst_req_1;
      W_ignq_2122_inst_ack_1<= rack(0);
      W_ignq_2122_inst : InterlockBuffer generic map ( -- 
        name => "W_ignq_2122_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => RPIPE_QUEUE_MONITOR_SIGNAL_2123_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ignq_2124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_2049_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2120_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2049_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2049_branch_req_0,
          ack0 => do_while_stmt_2049_branch_ack_0,
          ack1 => do_while_stmt_2049_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_2099_inst
    update_control_register_2100 <= (NOT_u1_u1_2095_wire and EQ_u8_u1_2098_wire);
    -- flow through binary operator AND_u1_u1_2106_inst
    set_globals_2107 <= (update_control_register_2100 and BITSEL_u32_u1_2105_wire);
    -- flow through binary operator BITSEL_u32_u1_2105_inst
    process(wdata_2075) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(wdata_2075, konst_2104_wire_constant, tmp_var);
      BITSEL_u32_u1_2105_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u33_2114_inst
    process(type_cast_2112_wire_constant, rdata_2091) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2112_wire_constant, rdata_2091, tmp_var);
      resp_2115 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_2098_inst
    process(index_2085) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_2085, konst_2097_wire_constant, tmp_var);
      EQ_u8_u1_2098_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2095_inst
    process(rwbar_2063) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rwbar_2063, tmp_var);
      NOT_u1_u1_2095_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_2052_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_2052_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_2052_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_2052_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_2052_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_2053 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- read from input-signal QUEUE_MONITOR_SIGNAL
    RPIPE_QUEUE_MONITOR_SIGNAL_2123_wire <= QUEUE_MONITOR_SIGNAL;
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_2116_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_2116_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_2116_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_2116_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_2116_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_2115;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_MAC_ENABLE_2029_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_MAC_ENABLE_2029_inst_req_0;
      WPIPE_MAC_ENABLE_2029_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_MAC_ENABLE_2029_inst_req_1;
      WPIPE_MAC_ENABLE_2029_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2030_wire_constant;
      MAC_ENABLE_write_1_gI: SplitGuardInterface generic map(name => "MAC_ENABLE_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      MAC_ENABLE_write_1: OutputPortRevised -- 
        generic map ( name => "MAC_ENABLE", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => MAC_ENABLE_pipe_write_req(0),
          oack => MAC_ENABLE_pipe_write_ack(0),
          odata => MAC_ENABLE_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_NIC_INTR_2032_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_INTR_2032_inst_req_0;
      WPIPE_NIC_INTR_2032_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_INTR_2032_inst_req_1;
      WPIPE_NIC_INTR_2032_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2033_wire_constant;
      NIC_INTR_write_2_gI: SplitGuardInterface generic map(name => "NIC_INTR_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_INTR_write_2: OutputPortRevised -- 
        generic map ( name => "NIC_INTR", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_INTR_pipe_write_req(0),
          oack => NIC_INTR_pipe_write_ack(0),
          odata => NIC_INTR_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_NIC_INTR_ENABLE_2035_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_INTR_ENABLE_2035_inst_req_0;
      WPIPE_NIC_INTR_ENABLE_2035_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_INTR_ENABLE_2035_inst_req_1;
      WPIPE_NIC_INTR_ENABLE_2035_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2036_wire_constant;
      NIC_INTR_ENABLE_write_3_gI: SplitGuardInterface generic map(name => "NIC_INTR_ENABLE_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_INTR_ENABLE_write_3: OutputPortRevised -- 
        generic map ( name => "NIC_INTR_ENABLE", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_INTR_ENABLE_pipe_write_req(0),
          oack => NIC_INTR_ENABLE_pipe_write_ack(0),
          odata => NIC_INTR_ENABLE_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_NIC_INTR_INTERNAL_2038_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_INTR_INTERNAL_2038_inst_req_0;
      WPIPE_NIC_INTR_INTERNAL_2038_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_INTR_INTERNAL_2038_inst_req_1;
      WPIPE_NIC_INTR_INTERNAL_2038_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2039_wire_constant;
      NIC_INTR_INTERNAL_write_4_gI: SplitGuardInterface generic map(name => "NIC_INTR_INTERNAL_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_INTR_INTERNAL_write_4: OutputPortRevised -- 
        generic map ( name => "NIC_INTR_INTERNAL", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_INTR_INTERNAL_pipe_write_req(0),
          oack => NIC_INTR_INTERNAL_pipe_write_ack(0),
          odata => NIC_INTR_INTERNAL_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_S_CONTROL_REGISTER_2041_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_S_CONTROL_REGISTER_2041_inst_req_0;
      WPIPE_S_CONTROL_REGISTER_2041_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_S_CONTROL_REGISTER_2041_inst_req_1;
      WPIPE_S_CONTROL_REGISTER_2041_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2042_wire_constant;
      S_CONTROL_REGISTER_write_5_gI: SplitGuardInterface generic map(name => "S_CONTROL_REGISTER_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      S_CONTROL_REGISTER_write_5: OutputPortRevised -- 
        generic map ( name => "S_CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => S_CONTROL_REGISTER_pipe_write_req(0),
          oack => S_CONTROL_REGISTER_pipe_write_ack(0),
          odata => S_CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_S_NUMBER_OF_SERVERS_2044_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_S_NUMBER_OF_SERVERS_2044_inst_req_0;
      WPIPE_S_NUMBER_OF_SERVERS_2044_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_S_NUMBER_OF_SERVERS_2044_inst_req_1;
      WPIPE_S_NUMBER_OF_SERVERS_2044_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2045_wire_constant;
      S_NUMBER_OF_SERVERS_write_6_gI: SplitGuardInterface generic map(name => "S_NUMBER_OF_SERVERS_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      S_NUMBER_OF_SERVERS_write_6: OutputPortRevised -- 
        generic map ( name => "S_NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => S_NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => S_NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => S_NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_memory_access_lock_2020_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_memory_access_lock_2020_inst_req_0;
      WPIPE_memory_access_lock_2020_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_memory_access_lock_2020_inst_req_1;
      WPIPE_memory_access_lock_2020_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2021_wire_constant;
      memory_access_lock_write_7_gI: SplitGuardInterface generic map(name => "memory_access_lock_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      memory_access_lock_write_7: OutputPortRevised -- 
        generic map ( name => "memory_access_lock", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => memory_access_lock_pipe_write_req(0),
          oack => memory_access_lock_pipe_write_ack(0),
          odata => memory_access_lock_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- shared call operator group (0) : call_stmt_2028_call 
    accessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(44 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2028_call_req_0;
      call_stmt_2028_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2028_call_req_1;
      call_stmt_2028_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_2023_wire_constant & konst_2024_wire_constant & konst_2025_wire_constant & konst_2026_wire_constant;
      ign_2028 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 45,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(1),
          ackR => accessRegister_call_acks(1),
          dataR => accessRegister_call_data(89 downto 45),
          tagR => accessRegister_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(1), -- cross-over
          ackL => accessRegister_return_reqs(1), -- cross-over
          dataL => accessRegister_return_data(63 downto 32),
          tagL => accessRegister_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2091_call 
    accessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(44 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2091_call_req_0;
      call_stmt_2091_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2091_call_req_1;
      call_stmt_2091_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rwbar_2063 & bmask_2067 & index_2085 & wdata_2075;
      rdata_2091 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 45,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2109_call 
    setGlobalSignals_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2109_call_req_0;
      call_stmt_2109_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2109_call_req_1;
      call_stmt_2109_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= set_globals_2107(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setGlobalSignals_call_group_2_gI: SplitGuardInterface generic map(name => "setGlobalSignals_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => setGlobalSignals_call_reqs(0),
          ackR => setGlobalSignals_call_acks(0),
          tagR => setGlobalSignals_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setGlobalSignals_return_acks(0), -- cross-over
          ackL => setGlobalSignals_return_reqs(0), -- cross-over
          tagL => setGlobalSignals_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end controlDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(9 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(9 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_2707_start: Boolean;
  signal delay_time_CP_2707_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1728_req_1 : boolean;
  signal do_while_stmt_1726_branch_ack_0 : boolean;
  signal T_1731_buf_req_1 : boolean;
  signal T_1731_buf_ack_1 : boolean;
  signal phi_stmt_1728_ack_0 : boolean;
  signal T_1731_buf_ack_0 : boolean;
  signal T_1731_buf_req_0 : boolean;
  signal phi_stmt_1728_req_0 : boolean;
  signal nR_1737_1730_buf_ack_1 : boolean;
  signal nR_1737_1730_buf_req_1 : boolean;
  signal nR_1737_1730_buf_ack_0 : boolean;
  signal nR_1737_1730_buf_req_0 : boolean;
  signal do_while_stmt_1726_branch_req_0 : boolean;
  signal do_while_stmt_1726_branch_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= delay_time_CP_2707_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  -- join of sample-req and update-req.. used to trigger CP.
  delay_time_CP_2707_start_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
    constant joinName: string(1 to 29) := "delay_time_CP_2707_start_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sample_req & update_req;
    gj_delay_time_CP_2707_start_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => delay_time_CP_2707_start, clk => clk, reset => reset); --
  end block;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_2707_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_2707: Block -- control-path 
    signal delay_time_CP_2707_elements: BooleanArray(34 downto 0);
    -- 
  begin -- 
    delay_time_CP_2707_elements(0) <= delay_time_CP_2707_start;
    delay_time_CP_2707_symbol <= delay_time_CP_2707_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1725/do_while_stmt_1726__entry__
      -- CP-element group 0: 	 branch_block_stmt_1725/branch_block_stmt_1725__entry__
      -- CP-element group 0: 	 branch_block_stmt_1725/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	34 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1725/do_while_stmt_1726__exit__
      -- CP-element group 1: 	 branch_block_stmt_1725/branch_block_stmt_1725__exit__
      -- CP-element group 1: 	 assign_stmt_1745/$exit
      -- CP-element group 1: 	 assign_stmt_1745/$entry
      -- CP-element group 1: 	 branch_block_stmt_1725/$exit
      -- CP-element group 1: 	 $exit
      -- 
    delay_time_CP_2707_elements(1) <= delay_time_CP_2707_elements(34);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726__entry__
      -- CP-element group 2: 	 branch_block_stmt_1725/do_while_stmt_1726/$entry
      -- 
    delay_time_CP_2707_elements(2) <= delay_time_CP_2707_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	34 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726__exit__
      -- 
    -- Element group delay_time_CP_2707_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_back
      -- 
    -- Element group delay_time_CP_2707_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	32 
    -- CP-element group 5: 	33 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1725/do_while_stmt_1726/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_taken/$entry
      -- 
    delay_time_CP_2707_elements(5) <= delay_time_CP_2707_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	31 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_body_done
      -- 
    delay_time_CP_2707_elements(6) <= delay_time_CP_2707_elements(31);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	17 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/back_edge_to_loop_body
      -- 
    delay_time_CP_2707_elements(7) <= delay_time_CP_2707_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	19 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/first_time_through_loop_body
      -- 
    delay_time_CP_2707_elements(8) <= delay_time_CP_2707_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	30 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/$entry
      -- 
    -- Element group delay_time_CP_2707_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	30 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/condition_evaluated
      -- 
    condition_evaluated_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(10), ack => do_while_stmt_1726_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2707_elements(16) & delay_time_CP_2707_elements(30);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2707_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_sample_req
      -- 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2707_elements(13) & delay_time_CP_2707_elements(16);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2707_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group delay_time_CP_2707_elements(12) is a control-delay.
    cp_element_12_delay: control_delay_element  generic map(name => " 12_delay", delay_value => 1)  port map(req => delay_time_CP_2707_elements(15), ack => delay_time_CP_2707_elements(12), clk => clk, reset =>reset);
    -- CP-element group 13:  join  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_start_
      -- 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2707_elements(9) & delay_time_CP_2707_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2707_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_start__ps
      -- CP-element group 14: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_update_req
      -- 
    delay_time_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2707_elements(9) & delay_time_CP_2707_elements(16);
      gj_delay_time_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2707_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_sample_ack
      -- 
    -- Element group delay_time_CP_2707_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/aggregated_phi_update_ack
      -- CP-element group 16: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_update_completed__ps
      -- 
    -- Element group delay_time_CP_2707_elements(16) is bound as output of CP function.
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	7 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_loopback_trigger
      -- 
    delay_time_CP_2707_elements(17) <= delay_time_CP_2707_elements(7);
    -- CP-element group 18:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_loopback_sample_req_ps
      -- CP-element group 18: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_loopback_sample_req
      -- 
    phi_stmt_1728_loopback_sample_req_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_loopback_sample_req_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(18), ack => phi_stmt_1728_req_0); -- 
    -- Element group delay_time_CP_2707_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_entry_trigger
      -- 
    delay_time_CP_2707_elements(19) <= delay_time_CP_2707_elements(8);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_entry_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_entry_sample_req_ps
      -- 
    phi_stmt_1728_entry_sample_req_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1728_entry_sample_req_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(20), ack => phi_stmt_1728_req_1); -- 
    -- Element group delay_time_CP_2707_elements(20) is bound as output of CP function.
    -- CP-element group 21:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_phi_mux_ack_ps
      -- CP-element group 21: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/phi_stmt_1728_phi_mux_ack
      -- 
    phi_stmt_1728_phi_mux_ack_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1728_ack_0, ack => delay_time_CP_2707_elements(21)); -- 
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Sample/req
      -- CP-element group 22: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_sample_start__ps
      -- 
    req_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(22), ack => nR_1737_1730_buf_req_0); -- 
    -- Element group delay_time_CP_2707_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Update/req
      -- CP-element group 23: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_update_start__ps
      -- 
    req_2771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(23), ack => nR_1737_1730_buf_req_1); -- 
    -- Element group delay_time_CP_2707_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Sample/ack
      -- CP-element group 24: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_sample_completed__ps
      -- 
    ack_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1737_1730_buf_ack_0, ack => delay_time_CP_2707_elements(24)); -- 
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Update/ack
      -- CP-element group 25: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_nR_1730_update_completed__ps
      -- 
    ack_2772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1737_1730_buf_ack_1, ack => delay_time_CP_2707_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Sample/req
      -- CP-element group 26: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_sample_start__ps
      -- 
    req_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(26), ack => T_1731_buf_req_0); -- 
    -- Element group delay_time_CP_2707_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Update/req
      -- CP-element group 27: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_update_start__ps
      -- 
    req_2789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2707_elements(27), ack => T_1731_buf_req_1); -- 
    -- Element group delay_time_CP_2707_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_sample_completed__ps
      -- 
    ack_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1731_buf_ack_0, ack => delay_time_CP_2707_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_Update/ack
      -- CP-element group 29: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/R_T_1731_update_completed__ps
      -- 
    ack_2790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1731_buf_ack_1, ack => delay_time_CP_2707_elements(29)); -- 
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	9 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	10 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group delay_time_CP_2707_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => delay_time_CP_2707_elements(9), ack => delay_time_CP_2707_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	6 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1725/do_while_stmt_1726/do_while_stmt_1726_loop_body/$exit
      -- 
    delay_time_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2707_elements(12) & delay_time_CP_2707_elements(15);
      gj_delay_time_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2707_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	5 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_exit/$exit
      -- CP-element group 32: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_exit/ack
      -- 
    ack_2796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1726_branch_ack_0, ack => delay_time_CP_2707_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	5 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_taken/$exit
      -- CP-element group 33: 	 branch_block_stmt_1725/do_while_stmt_1726/loop_taken/ack
      -- 
    ack_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1726_branch_ack_1, ack => delay_time_CP_2707_elements(33)); -- 
    -- CP-element group 34:  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	3 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	1 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1725/do_while_stmt_1726/$exit
      -- 
    delay_time_CP_2707_elements(34) <= delay_time_CP_2707_elements(3);
    delay_time_do_while_stmt_1726_terminator_2801: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_1726_terminator_2801", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_2707_elements(6),loop_continue => delay_time_CP_2707_elements(33),loop_terminate => delay_time_CP_2707_elements(32),loop_back => delay_time_CP_2707_elements(4),loop_exit => delay_time_CP_2707_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1728_phi_seq_2791_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_2707_elements(17);
      delay_time_CP_2707_elements(22)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_2707_elements(24);
      delay_time_CP_2707_elements(23)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_2707_elements(25);
      delay_time_CP_2707_elements(18) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_2707_elements(19);
      delay_time_CP_2707_elements(26)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_2707_elements(28);
      delay_time_CP_2707_elements(27)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_2707_elements(29);
      delay_time_CP_2707_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1728_phi_seq_2791 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1728_phi_seq_2791") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_2707_elements(11), 
          phi_sample_ack => delay_time_CP_2707_elements(15), 
          phi_update_req => delay_time_CP_2707_elements(14), 
          phi_update_ack => delay_time_CP_2707_elements(16), 
          phi_mux_ack => delay_time_CP_2707_elements(21), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2732_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_2707_elements(7);
        preds(1)  <= delay_time_CP_2707_elements(8);
        entry_tmerge_2732 : transition_merge -- 
          generic map(name => " entry_tmerge_2732")
          port map (preds => preds, symbol_out => delay_time_CP_2707_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_1728 : std_logic_vector(9 downto 0);
    signal T_1731_buffered : std_logic_vector(9 downto 0);
    signal UGT_u10_u1_1741_wire : std_logic_vector(0 downto 0);
    signal konst_1735_wire_constant : std_logic_vector(9 downto 0);
    signal konst_1740_wire_constant : std_logic_vector(9 downto 0);
    signal nR_1737 : std_logic_vector(9 downto 0);
    signal nR_1737_1730_buffered : std_logic_vector(9 downto 0);
    -- 
  begin -- 
    konst_1735_wire_constant <= "0000000001";
    konst_1740_wire_constant <= "0000000000";
    phi_stmt_1728: Block -- phi operator 
      signal idata: std_logic_vector(19 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nR_1737_1730_buffered & T_1731_buffered;
      req <= phi_stmt_1728_req_0 & phi_stmt_1728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1728",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 10) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1728_ack_0,
          idata => idata,
          odata => R_1728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1728
    T_1731_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_1731_buf_req_0;
      T_1731_buf_ack_0<= wack(0);
      rreq(0) <= T_1731_buf_req_1;
      T_1731_buf_ack_1<= rack(0);
      T_1731_buf : InterlockBuffer generic map ( -- 
        name => "T_1731_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 10,
        out_data_width => 10,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_1731_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nR_1737_1730_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_1737_1730_buf_req_0;
      nR_1737_1730_buf_ack_0<= wack(0);
      rreq(0) <= nR_1737_1730_buf_req_1;
      nR_1737_1730_buf_ack_1<= rack(0);
      nR_1737_1730_buf : InterlockBuffer generic map ( -- 
        name => "nR_1737_1730_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 10,
        out_data_width => 10,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_1737,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_1737_1730_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1726_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u10_u1_1741_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1726_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1726_branch_req_0,
          ack0 => do_while_stmt_1726_branch_ack_0,
          ack1 => do_while_stmt_1726_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator SUB_u10_u10_1736_inst
    nR_1737 <= std_logic_vector(unsigned(R_1728) - unsigned(konst_1735_wire_constant));
    -- flow through binary operator UGT_u10_u1_1741_inst
    process(R_1728) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_1728, konst_1740_wire_constant, tmp_var);
      UGT_u10_u1_1741_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity doMemAccess is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    opcode : in  std_logic_vector(2 downto 0);
    base_addr : in  std_logic_vector(63 downto 0);
    offset : in  std_logic_vector(63 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    memory_access_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
    memory_access_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
    memory_access_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
    memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
    memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
    memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
    accessMemoryWordBase_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWordBase_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWordBase_call_data : out  std_logic_vector(169 downto 0);
    accessMemoryWordBase_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWordBase_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWordBase_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWordBase_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWordBase_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemoryByteBase_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryByteBase_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryByteBase_call_data : out  std_logic_vector(145 downto 0);
    accessMemoryByteBase_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemoryByteBase_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryByteBase_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryByteBase_return_data : in   std_logic_vector(7 downto 0);
    accessMemoryByteBase_return_tag :  in   std_logic_vector(1 downto 0);
    accessMemoryDwordBase_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDwordBase_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDwordBase_call_data : out  std_logic_vector(201 downto 0);
    accessMemoryDwordBase_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryDwordBase_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDwordBase_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDwordBase_return_data : in   std_logic_vector(63 downto 0);
    accessMemoryDwordBase_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity doMemAccess;
architecture doMemAccess_arch of doMemAccess is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 203)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal opcode_buffer :  std_logic_vector(2 downto 0);
  signal opcode_update_enable: Boolean;
  signal base_addr_buffer :  std_logic_vector(63 downto 0);
  signal base_addr_update_enable: Boolean;
  signal offset_buffer :  std_logic_vector(63 downto 0);
  signal offset_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal doMemAccess_CP_742_start: Boolean;
  signal doMemAccess_CP_742_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryWordBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
      calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
      calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
      calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
      accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
      accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryByteBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      byte_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wbyte : in  std_logic_vector(7 downto 0);
      rbyte : out  std_logic_vector(7 downto 0);
      calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
      calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
      calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
      calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
      accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
      accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryDwordBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
      calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
      calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
      calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
      accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
      accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_base_addr_716_delayed_17_0_766_inst_req_0 : boolean;
  signal W_base_addr_716_delayed_17_0_766_inst_ack_1 : boolean;
  signal call_stmt_749_call_req_0 : boolean;
  signal W_is_ldstub_709_delayed_17_0_760_inst_req_1 : boolean;
  signal call_stmt_749_call_req_1 : boolean;
  signal W_base_addr_716_delayed_17_0_766_inst_ack_0 : boolean;
  signal RPIPE_memory_access_lock_706_inst_req_0 : boolean;
  signal call_stmt_749_call_ack_1 : boolean;
  signal W_is_ldstub_664_delayed_1_0_709_inst_req_1 : boolean;
  signal call_stmt_737_call_req_1 : boolean;
  signal RPIPE_memory_access_lock_706_inst_ack_0 : boolean;
  signal call_stmt_725_call_req_0 : boolean;
  signal call_stmt_737_call_ack_1 : boolean;
  signal RPIPE_memory_access_lock_706_inst_req_1 : boolean;
  signal W_offset_717_delayed_17_0_769_inst_ack_1 : boolean;
  signal W_tag_710_delayed_17_0_763_inst_req_1 : boolean;
  signal W_tag_710_delayed_17_0_763_inst_ack_1 : boolean;
  signal W_is_ldstub_703_delayed_17_0_750_inst_ack_0 : boolean;
  signal W_is_ldstub_703_delayed_17_0_750_inst_req_1 : boolean;
  signal call_stmt_725_call_ack_1 : boolean;
  signal OR_u1_u1_787_inst_req_0 : boolean;
  signal W_is_ldstub_703_delayed_17_0_750_inst_ack_1 : boolean;
  signal W_is_ldstub_664_delayed_1_0_709_inst_ack_1 : boolean;
  signal W_tag_710_delayed_17_0_763_inst_req_0 : boolean;
  signal W_is_ldstub_709_delayed_17_0_760_inst_ack_0 : boolean;
  signal W_is_ldstub_709_delayed_17_0_760_inst_req_0 : boolean;
  signal W_is_ldstub_709_delayed_17_0_760_inst_ack_1 : boolean;
  signal W_base_addr_716_delayed_17_0_766_inst_req_1 : boolean;
  signal call_stmt_725_call_ack_0 : boolean;
  signal W_tag_710_delayed_17_0_763_inst_ack_0 : boolean;
  signal call_stmt_737_call_req_0 : boolean;
  signal call_stmt_725_call_req_1 : boolean;
  signal W_offset_717_delayed_17_0_769_inst_req_1 : boolean;
  signal WPIPE_memory_access_lock_713_inst_ack_1 : boolean;
  signal W_offset_717_delayed_17_0_769_inst_req_0 : boolean;
  signal W_is_ldstub_664_delayed_1_0_709_inst_ack_0 : boolean;
  signal WPIPE_memory_access_lock_713_inst_req_1 : boolean;
  signal RPIPE_memory_access_lock_706_inst_ack_1 : boolean;
  signal W_is_ldstub_664_delayed_1_0_709_inst_req_0 : boolean;
  signal WPIPE_memory_access_lock_713_inst_ack_0 : boolean;
  signal W_offset_717_delayed_17_0_769_inst_ack_0 : boolean;
  signal call_stmt_749_call_ack_0 : boolean;
  signal WPIPE_memory_access_lock_713_inst_req_0 : boolean;
  signal W_is_ldstub_703_delayed_17_0_750_inst_req_0 : boolean;
  signal call_stmt_783_call_req_0 : boolean;
  signal call_stmt_783_call_ack_0 : boolean;
  signal call_stmt_783_call_req_1 : boolean;
  signal call_stmt_783_call_ack_1 : boolean;
  signal call_stmt_737_call_ack_0 : boolean;
  signal OR_u1_u1_787_inst_ack_0 : boolean;
  signal OR_u1_u1_787_inst_req_1 : boolean;
  signal OR_u1_u1_787_inst_ack_1 : boolean;
  signal W_is_word_access_731_delayed_17_0_789_inst_req_0 : boolean;
  signal W_is_word_access_731_delayed_17_0_789_inst_ack_0 : boolean;
  signal W_is_word_access_731_delayed_17_0_789_inst_req_1 : boolean;
  signal W_is_word_access_731_delayed_17_0_789_inst_ack_1 : boolean;
  signal W_is_dword_access_739_delayed_16_0_792_inst_req_0 : boolean;
  signal W_is_dword_access_739_delayed_16_0_792_inst_ack_0 : boolean;
  signal W_is_dword_access_739_delayed_16_0_792_inst_req_1 : boolean;
  signal W_is_dword_access_739_delayed_16_0_792_inst_ack_1 : boolean;
  signal MUX_799_inst_req_0 : boolean;
  signal MUX_799_inst_ack_0 : boolean;
  signal MUX_799_inst_req_1 : boolean;
  signal MUX_799_inst_ack_1 : boolean;
  signal WPIPE_memory_access_lock_822_inst_req_0 : boolean;
  signal WPIPE_memory_access_lock_822_inst_ack_0 : boolean;
  signal WPIPE_memory_access_lock_822_inst_req_1 : boolean;
  signal WPIPE_memory_access_lock_822_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "doMemAccess_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 203) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(10 downto 8) <= opcode;
  opcode_buffer <= in_buffer_data_out(10 downto 8);
  in_buffer_data_in(74 downto 11) <= base_addr;
  base_addr_buffer <= in_buffer_data_out(74 downto 11);
  in_buffer_data_in(138 downto 75) <= offset;
  offset_buffer <= in_buffer_data_out(138 downto 75);
  in_buffer_data_in(202 downto 139) <= wdata;
  wdata_buffer <= in_buffer_data_out(202 downto 139);
  in_buffer_data_in(tag_length + 202 downto 203) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 202 downto 203);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= tag_update_enable & opcode_update_enable & base_addr_update_enable & offset_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  doMemAccess_CP_742_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "doMemAccess_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= doMemAccess_CP_742_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= doMemAccess_CP_742_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= doMemAccess_CP_742_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  doMemAccess_CP_742: Block -- control-path 
    signal doMemAccess_CP_742_elements: BooleanArray(82 downto 0);
    -- 
  begin -- 
    doMemAccess_CP_742_elements(0) <= doMemAccess_CP_742_start;
    doMemAccess_CP_742_symbol <= doMemAccess_CP_742_elements(82);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	28 
    -- CP-element group 1: 	32 
    -- CP-element group 1: 	36 
    -- CP-element group 1: 	12 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	40 
    -- CP-element group 1: 	44 
    -- CP-element group 1: 	48 
    -- CP-element group 1: 	56 
    -- CP-element group 1: 	60 
    -- CP-element group 1: 	64 
    -- CP-element group 1: 	73 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_640_to_assign_stmt_825/$entry
      -- 
    doMemAccess_CP_742_elements(1) <= doMemAccess_CP_742_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	42 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	76 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_825/tag_update_enable
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_825/tag_update_enable_out
      -- 
    doMemAccess_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(22) & doMemAccess_CP_742_elements(26) & doMemAccess_CP_742_elements(30) & doMemAccess_CP_742_elements(42);
      gj_doMemAccess_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	22 
    -- CP-element group 3: 	26 
    -- CP-element group 3: 	30 
    -- CP-element group 3: 	34 
    -- CP-element group 3: 	14 
    -- CP-element group 3: 	38 
    -- CP-element group 3: 	58 
    -- CP-element group 3: 	62 
    -- CP-element group 3: 	66 
    -- CP-element group 3: 	74 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	77 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_640_to_assign_stmt_825/opcode_update_enable
      -- CP-element group 3: 	 assign_stmt_640_to_assign_stmt_825/opcode_update_enable_out
      -- 
    doMemAccess_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(22) & doMemAccess_CP_742_elements(26) & doMemAccess_CP_742_elements(30) & doMemAccess_CP_742_elements(34) & doMemAccess_CP_742_elements(14) & doMemAccess_CP_742_elements(38) & doMemAccess_CP_742_elements(58) & doMemAccess_CP_742_elements(62) & doMemAccess_CP_742_elements(66) & doMemAccess_CP_742_elements(74);
      gj_doMemAccess_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	22 
    -- CP-element group 4: 	26 
    -- CP-element group 4: 	30 
    -- CP-element group 4: 	46 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	78 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_640_to_assign_stmt_825/base_addr_update_enable_out
      -- CP-element group 4: 	 assign_stmt_640_to_assign_stmt_825/base_addr_update_enable
      -- 
    doMemAccess_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(22) & doMemAccess_CP_742_elements(26) & doMemAccess_CP_742_elements(30) & doMemAccess_CP_742_elements(46);
      gj_doMemAccess_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	22 
    -- CP-element group 5: 	26 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	50 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	79 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_640_to_assign_stmt_825/offset_update_enable_out
      -- CP-element group 5: 	 assign_stmt_640_to_assign_stmt_825/offset_update_enable
      -- 
    doMemAccess_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(22) & doMemAccess_CP_742_elements(26) & doMemAccess_CP_742_elements(30) & doMemAccess_CP_742_elements(50);
      gj_doMemAccess_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	22 
    -- CP-element group 6: 	26 
    -- CP-element group 6: 	30 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	80 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_640_to_assign_stmt_825/wdata_update_enable
      -- CP-element group 6: 	 assign_stmt_640_to_assign_stmt_825/wdata_update_enable_out
      -- 
    doMemAccess_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(22) & doMemAccess_CP_742_elements(26) & doMemAccess_CP_742_elements(30);
      gj_doMemAccess_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	81 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	25 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	69 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_640_to_assign_stmt_825/rdata_update_enable
      -- CP-element group 7: 	 assign_stmt_640_to_assign_stmt_825/rdata_update_enable_in
      -- 
    doMemAccess_CP_742_elements(7) <= doMemAccess_CP_742_elements(81);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	11 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Sample/rr
      -- CP-element group 8: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_sample_start_
      -- CP-element group 8: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Sample/$entry
      -- 
    rr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(8), ack => RPIPE_memory_access_lock_706_inst_req_0); -- 
    doMemAccess_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(11);
      gj_doMemAccess_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	17 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_update_start_
      -- CP-element group 9: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Update/cr
      -- CP-element group 9: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Update/$entry
      -- 
    cr_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(9), ack => RPIPE_memory_access_lock_706_inst_req_1); -- 
    doMemAccess_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "doMemAccess_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(10) & doMemAccess_CP_742_elements(17);
      gj_doMemAccess_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	9 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_sample_completed_
      -- CP-element group 10: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Sample/ra
      -- CP-element group 10: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Sample/$exit
      -- 
    ra_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_memory_access_lock_706_inst_ack_0, ack => doMemAccess_CP_742_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	8 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_update_completed_
      -- CP-element group 11: 	 assign_stmt_640_to_assign_stmt_825/barrier_stmt_708_update_completed_
      -- CP-element group 11: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Update/$exit
      -- CP-element group 11: 	 assign_stmt_640_to_assign_stmt_825/RPIPE_memory_access_lock_706_Update/ca
      -- 
    ca_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_memory_access_lock_706_inst_ack_1, ack => doMemAccess_CP_742_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: 	1 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Sample/req
      -- CP-element group 12: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Sample/$entry
      -- CP-element group 12: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_sample_start_
      -- 
    req_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(12), ack => W_is_ldstub_664_delayed_1_0_709_inst_req_0); -- 
    doMemAccess_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(11) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(14);
      gj_doMemAccess_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Update/req
      -- CP-element group 13: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Update/$entry
      -- CP-element group 13: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_update_start_
      -- 
    req_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(13), ack => W_is_ldstub_664_delayed_1_0_709_inst_req_1); -- 
    doMemAccess_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(15) & doMemAccess_CP_742_elements(17);
      gj_doMemAccess_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_sample_completed_
      -- CP-element group 14: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Sample/ack
      -- CP-element group 14: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Sample/$exit
      -- 
    ack_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_ldstub_664_delayed_1_0_709_inst_ack_0, ack => doMemAccess_CP_742_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	19 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Update/$exit
      -- CP-element group 15: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_Update/ack
      -- CP-element group 15: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_711_update_completed_
      -- 
    ack_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_ldstub_664_delayed_1_0_709_inst_ack_1, ack => doMemAccess_CP_742_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: 	11 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	75 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_sample_start_
      -- CP-element group 16: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Sample/req
      -- 
    req_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(16), ack => WPIPE_memory_access_lock_713_inst_req_0); -- 
    doMemAccess_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(15) & doMemAccess_CP_742_elements(11) & doMemAccess_CP_742_elements(18) & doMemAccess_CP_742_elements(75);
      gj_doMemAccess_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17: 	9 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_update_start_
      -- CP-element group 17: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_sample_completed_
      -- CP-element group 17: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Sample/$exit
      -- CP-element group 17: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Update/req
      -- CP-element group 17: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Update/$entry
      -- CP-element group 17: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Sample/ack
      -- 
    ack_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_memory_access_lock_713_inst_ack_0, ack => doMemAccess_CP_742_elements(17)); -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(17), ack => WPIPE_memory_access_lock_713_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	73 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_update_completed_
      -- CP-element group 18: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Update/ack
      -- CP-element group 18: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_713_Update/$exit
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_memory_access_lock_713_inst_ack_1, ack => doMemAccess_CP_742_elements(18)); -- 
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	32 
    -- CP-element group 19: 	36 
    -- CP-element group 19: 	40 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	48 
    -- CP-element group 19: 	56 
    -- CP-element group 19: 	60 
    -- CP-element group 19: 	64 
    -- CP-element group 19: 	68 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 assign_stmt_640_to_assign_stmt_825/barrier_stmt_716_update_completed_
      -- 
    doMemAccess_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(15) & doMemAccess_CP_742_elements(18);
      gj_doMemAccess_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	1 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: 	55 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Sample/crr
      -- CP-element group 20: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Sample/$entry
      -- CP-element group 20: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_sample_start_
      -- 
    crr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(20), ack => call_stmt_725_call_req_0); -- 
    doMemAccess_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(22) & doMemAccess_CP_742_elements(55);
      gj_doMemAccess_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	54 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Update/ccr
      -- CP-element group 21: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_update_start_
      -- CP-element group 21: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Update/$entry
      -- 
    ccr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(21), ack => call_stmt_725_call_req_1); -- 
    doMemAccess_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(7) & doMemAccess_CP_742_elements(23) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	4 
    -- CP-element group 22: 	2 
    -- CP-element group 22: 	5 
    -- CP-element group 22: 	6 
    -- CP-element group 22: 	3 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Sample/$exit
      -- CP-element group 22: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Sample/cra
      -- CP-element group 22: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_sample_completed_
      -- 
    cra_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_725_call_ack_0, ack => doMemAccess_CP_742_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	52 
    -- CP-element group 23: 	72 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Update/cca
      -- CP-element group 23: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_update_completed_
      -- CP-element group 23: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_725_Update/$exit
      -- 
    cca_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_725_call_ack_1, ack => doMemAccess_CP_742_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Sample/$entry
      -- CP-element group 24: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Sample/crr
      -- CP-element group 24: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_sample_start_
      -- 
    crr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(24), ack => call_stmt_737_call_req_0); -- 
    doMemAccess_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(23) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(26);
      gj_doMemAccess_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	7 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Update/ccr
      -- CP-element group 25: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Update/$entry
      -- CP-element group 25: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_update_start_
      -- 
    ccr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(25), ack => call_stmt_737_call_req_1); -- 
    doMemAccess_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(7) & doMemAccess_CP_742_elements(27);
      gj_doMemAccess_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	4 
    -- CP-element group 26: 	2 
    -- CP-element group 26: 	5 
    -- CP-element group 26: 	6 
    -- CP-element group 26: 	3 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Sample/$exit
      -- CP-element group 26: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_sample_completed_
      -- CP-element group 26: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Sample/cra
      -- 
    cra_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_737_call_ack_0, ack => doMemAccess_CP_742_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	72 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Update/cca
      -- CP-element group 27: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_Update/$exit
      -- CP-element group 27: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_737_update_completed_
      -- 
    cca_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_737_call_ack_1, ack => doMemAccess_CP_742_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: 	1 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Sample/crr
      -- CP-element group 28: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_sample_start_
      -- CP-element group 28: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Sample/$entry
      -- 
    crr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(28), ack => call_stmt_749_call_req_0); -- 
    doMemAccess_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(27) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(30);
      gj_doMemAccess_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: 	70 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Update/ccr
      -- CP-element group 29: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Update/$entry
      -- CP-element group 29: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_update_start_
      -- 
    ccr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(29), ack => call_stmt_749_call_req_1); -- 
    doMemAccess_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(31) & doMemAccess_CP_742_elements(70);
      gj_doMemAccess_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: 	4 
    -- CP-element group 30: 	2 
    -- CP-element group 30: 	5 
    -- CP-element group 30: 	6 
    -- CP-element group 30: 	3 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Sample/$exit
      -- CP-element group 30: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Sample/cra
      -- CP-element group 30: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_sample_completed_
      -- 
    cra_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_749_call_ack_0, ack => doMemAccess_CP_742_elements(30)); -- 
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	52 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	72 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Update/cca
      -- CP-element group 31: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_Update/$exit
      -- CP-element group 31: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_749_update_completed_
      -- 
    cca_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_749_call_ack_1, ack => doMemAccess_CP_742_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	19 
    -- CP-element group 32: 	1 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Sample/req
      -- CP-element group 32: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Sample/$entry
      -- CP-element group 32: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_sample_start_
      -- 
    req_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(32), ack => W_is_ldstub_703_delayed_17_0_750_inst_req_0); -- 
    doMemAccess_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(34);
      gj_doMemAccess_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: 	54 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Update/$entry
      -- CP-element group 33: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Update/req
      -- CP-element group 33: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_update_start_
      -- 
    req_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(33), ack => W_is_ldstub_703_delayed_17_0_750_inst_req_1); -- 
    doMemAccess_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(35) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: 	3 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Sample/ack
      -- CP-element group 34: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Sample/$exit
      -- CP-element group 34: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_sample_completed_
      -- 
    ack_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_ldstub_703_delayed_17_0_750_inst_ack_0, ack => doMemAccess_CP_742_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	52 
    -- CP-element group 35: 	72 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Update/$exit
      -- CP-element group 35: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_update_completed_
      -- CP-element group 35: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_752_Update/ack
      -- 
    ack_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_ldstub_703_delayed_17_0_750_inst_ack_1, ack => doMemAccess_CP_742_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	19 
    -- CP-element group 36: 	1 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_sample_start_
      -- CP-element group 36: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Sample/req
      -- 
    req_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(36), ack => W_is_ldstub_709_delayed_17_0_760_inst_req_0); -- 
    doMemAccess_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(38);
      gj_doMemAccess_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Update/req
      -- CP-element group 37: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_update_start_
      -- CP-element group 37: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Update/$entry
      -- 
    req_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(37), ack => W_is_ldstub_709_delayed_17_0_760_inst_req_1); -- 
    doMemAccess_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(39) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: 	3 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_sample_completed_
      -- CP-element group 38: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Sample/ack
      -- 
    ack_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_ldstub_709_delayed_17_0_760_inst_ack_0, ack => doMemAccess_CP_742_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: 	72 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_update_completed_
      -- CP-element group 39: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Update/ack
      -- CP-element group 39: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_762_Update/$exit
      -- 
    ack_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_ldstub_709_delayed_17_0_760_inst_ack_1, ack => doMemAccess_CP_742_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	19 
    -- CP-element group 40: 	1 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Sample/req
      -- CP-element group 40: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_sample_start_
      -- 
    req_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(40), ack => W_tag_710_delayed_17_0_763_inst_req_0); -- 
    doMemAccess_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(42);
      gj_doMemAccess_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	54 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Update/$entry
      -- CP-element group 41: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Update/req
      -- CP-element group 41: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_update_start_
      -- 
    req_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(41), ack => W_tag_710_delayed_17_0_763_inst_req_1); -- 
    doMemAccess_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(43) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	2 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Sample/ack
      -- CP-element group 42: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_sample_completed_
      -- 
    ack_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_710_delayed_17_0_763_inst_ack_0, ack => doMemAccess_CP_742_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	52 
    -- CP-element group 43: 	72 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Update/$exit
      -- CP-element group 43: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_Update/ack
      -- CP-element group 43: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_765_update_completed_
      -- 
    ack_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_710_delayed_17_0_763_inst_ack_1, ack => doMemAccess_CP_742_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	19 
    -- CP-element group 44: 	1 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Sample/req
      -- CP-element group 44: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_sample_start_
      -- CP-element group 44: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Sample/$entry
      -- 
    req_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(44), ack => W_base_addr_716_delayed_17_0_766_inst_req_0); -- 
    doMemAccess_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(46);
      gj_doMemAccess_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	54 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_update_start_
      -- CP-element group 45: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Update/req
      -- CP-element group 45: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Update/$entry
      -- 
    req_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(45), ack => W_base_addr_716_delayed_17_0_766_inst_req_1); -- 
    doMemAccess_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(47) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	4 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Sample/ack
      -- CP-element group 46: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_sample_completed_
      -- 
    ack_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_addr_716_delayed_17_0_766_inst_ack_0, ack => doMemAccess_CP_742_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	52 
    -- CP-element group 47: 	72 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Update/ack
      -- CP-element group 47: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_Update/$exit
      -- CP-element group 47: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_768_update_completed_
      -- 
    ack_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_addr_716_delayed_17_0_766_inst_ack_1, ack => doMemAccess_CP_742_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	19 
    -- CP-element group 48: 	1 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_sample_start_
      -- CP-element group 48: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Sample/req
      -- CP-element group 48: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Sample/$entry
      -- 
    req_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(48), ack => W_offset_717_delayed_17_0_769_inst_req_0); -- 
    doMemAccess_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(50);
      gj_doMemAccess_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	54 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Update/$entry
      -- CP-element group 49: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_update_start_
      -- CP-element group 49: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Update/req
      -- 
    req_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(49), ack => W_offset_717_delayed_17_0_769_inst_req_1); -- 
    doMemAccess_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(51) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_sample_completed_
      -- CP-element group 50: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Sample/ack
      -- 
    ack_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_offset_717_delayed_17_0_769_inst_ack_0, ack => doMemAccess_CP_742_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	72 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Update/ack
      -- CP-element group 51: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_update_completed_
      -- CP-element group 51: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_771_Update/$exit
      -- 
    ack_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_offset_717_delayed_17_0_769_inst_ack_1, ack => doMemAccess_CP_742_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	23 
    -- CP-element group 52: 	31 
    -- CP-element group 52: 	35 
    -- CP-element group 52: 	39 
    -- CP-element group 52: 	43 
    -- CP-element group 52: 	47 
    -- CP-element group 52: 	51 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_sample_start_
      -- CP-element group 52: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Sample/crr
      -- CP-element group 52: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Sample/$entry
      -- 
    crr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(52), ack => call_stmt_783_call_req_0); -- 
    doMemAccess_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(23) & doMemAccess_CP_742_elements(31) & doMemAccess_CP_742_elements(35) & doMemAccess_CP_742_elements(39) & doMemAccess_CP_742_elements(43) & doMemAccess_CP_742_elements(47) & doMemAccess_CP_742_elements(51) & doMemAccess_CP_742_elements(54);
      gj_doMemAccess_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Update/ccr
      -- CP-element group 53: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Update/$entry
      -- CP-element group 53: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_update_start_
      -- 
    ccr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(53), ack => call_stmt_783_call_req_1); -- 
    doMemAccess_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= doMemAccess_CP_742_elements(55);
      gj_doMemAccess_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	21 
    -- CP-element group 54: 	33 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	41 
    -- CP-element group 54: 	45 
    -- CP-element group 54: 	49 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_sample_completed_
      -- CP-element group 54: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Sample/cra
      -- CP-element group 54: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Sample/$exit
      -- 
    cra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_783_call_ack_0, ack => doMemAccess_CP_742_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	72 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	20 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Update/$exit
      -- CP-element group 55: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_update_completed_
      -- CP-element group 55: 	 assign_stmt_640_to_assign_stmt_825/call_stmt_783_Update/cca
      -- 
    cca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_783_call_ack_1, ack => doMemAccess_CP_742_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	19 
    -- CP-element group 56: 	1 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Sample/rr
      -- CP-element group 56: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_sample_start_
      -- 
    rr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(56), ack => OR_u1_u1_787_inst_req_0); -- 
    doMemAccess_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(58);
      gj_doMemAccess_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_update_start_
      -- CP-element group 57: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Update/$entry
      -- CP-element group 57: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Update/cr
      -- 
    cr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(57), ack => OR_u1_u1_787_inst_req_1); -- 
    doMemAccess_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(7) & doMemAccess_CP_742_elements(59);
      gj_doMemAccess_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	3 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Sample/$exit
      -- CP-element group 58: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_sample_completed_
      -- CP-element group 58: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Sample/ra
      -- 
    ra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_787_inst_ack_0, ack => doMemAccess_CP_742_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	72 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_update_completed_
      -- CP-element group 59: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Update/$exit
      -- CP-element group 59: 	 assign_stmt_640_to_assign_stmt_825/OR_u1_u1_787_Update/ca
      -- 
    ca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_787_inst_ack_1, ack => doMemAccess_CP_742_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	19 
    -- CP-element group 60: 	1 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_sample_start_
      -- CP-element group 60: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Sample/$entry
      -- CP-element group 60: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Sample/req
      -- 
    req_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(60), ack => W_is_word_access_731_delayed_17_0_789_inst_req_0); -- 
    doMemAccess_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(62);
      gj_doMemAccess_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_update_start_
      -- CP-element group 61: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Update/$entry
      -- CP-element group 61: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Update/req
      -- 
    req_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(61), ack => W_is_word_access_731_delayed_17_0_789_inst_req_1); -- 
    doMemAccess_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(7) & doMemAccess_CP_742_elements(63);
      gj_doMemAccess_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	3 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_sample_completed_
      -- CP-element group 62: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Sample/ack
      -- 
    ack_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_word_access_731_delayed_17_0_789_inst_ack_0, ack => doMemAccess_CP_742_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	72 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_update_completed_
      -- CP-element group 63: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Update/$exit
      -- CP-element group 63: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_791_Update/ack
      -- 
    ack_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_word_access_731_delayed_17_0_789_inst_ack_1, ack => doMemAccess_CP_742_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	19 
    -- CP-element group 64: 	1 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_sample_start_
      -- CP-element group 64: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Sample/req
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(64), ack => W_is_dword_access_739_delayed_16_0_792_inst_req_0); -- 
    doMemAccess_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(66);
      gj_doMemAccess_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	70 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_update_start_
      -- CP-element group 65: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Update/$entry
      -- CP-element group 65: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Update/req
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(65), ack => W_is_dword_access_739_delayed_16_0_792_inst_req_1); -- 
    doMemAccess_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(67) & doMemAccess_CP_742_elements(70);
      gj_doMemAccess_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_sample_completed_
      -- CP-element group 66: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Sample/ack
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_dword_access_739_delayed_16_0_792_inst_ack_0, ack => doMemAccess_CP_742_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	72 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_update_completed_
      -- CP-element group 67: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Update/$exit
      -- CP-element group 67: 	 assign_stmt_640_to_assign_stmt_825/assign_stmt_794_Update/ack
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_is_dword_access_739_delayed_16_0_792_inst_ack_1, ack => doMemAccess_CP_742_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	19 
    -- CP-element group 68: 	31 
    -- CP-element group 68: 	67 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_sample_start_
      -- CP-element group 68: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_start/$entry
      -- CP-element group 68: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_start/req
      -- 
    req_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(68), ack => MUX_799_inst_req_0); -- 
    doMemAccess_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(19) & doMemAccess_CP_742_elements(31) & doMemAccess_CP_742_elements(67) & doMemAccess_CP_742_elements(70);
      gj_doMemAccess_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	7 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_update_start_
      -- CP-element group 69: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_complete/$entry
      -- CP-element group 69: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_complete/req
      -- 
    req_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(69), ack => MUX_799_inst_req_1); -- 
    doMemAccess_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(7) & doMemAccess_CP_742_elements(71);
      gj_doMemAccess_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_sample_completed_
      -- CP-element group 70: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_start/$exit
      -- CP-element group 70: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_start/ack
      -- 
    ack_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_799_inst_ack_0, ack => doMemAccess_CP_742_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_update_completed_
      -- CP-element group 71: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_complete/$exit
      -- CP-element group 71: 	 assign_stmt_640_to_assign_stmt_825/MUX_799_complete/ack
      -- 
    ack_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_799_inst_ack_1, ack => doMemAccess_CP_742_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	23 
    -- CP-element group 72: 	27 
    -- CP-element group 72: 	31 
    -- CP-element group 72: 	35 
    -- CP-element group 72: 	39 
    -- CP-element group 72: 	43 
    -- CP-element group 72: 	47 
    -- CP-element group 72: 	51 
    -- CP-element group 72: 	55 
    -- CP-element group 72: 	59 
    -- CP-element group 72: 	63 
    -- CP-element group 72: 	67 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 assign_stmt_640_to_assign_stmt_825/barrier_stmt_820_update_completed_
      -- 
    doMemAccess_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 15,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(23) & doMemAccess_CP_742_elements(27) & doMemAccess_CP_742_elements(31) & doMemAccess_CP_742_elements(35) & doMemAccess_CP_742_elements(39) & doMemAccess_CP_742_elements(43) & doMemAccess_CP_742_elements(47) & doMemAccess_CP_742_elements(51) & doMemAccess_CP_742_elements(55) & doMemAccess_CP_742_elements(59) & doMemAccess_CP_742_elements(63) & doMemAccess_CP_742_elements(67) & doMemAccess_CP_742_elements(71);
      gj_doMemAccess_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	18 
    -- CP-element group 73: 	1 
    -- CP-element group 73: 	72 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_sample_start_
      -- CP-element group 73: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Sample/$entry
      -- CP-element group 73: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Sample/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(73), ack => WPIPE_memory_access_lock_822_inst_req_0); -- 
    doMemAccess_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "doMemAccess_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= doMemAccess_CP_742_elements(18) & doMemAccess_CP_742_elements(1) & doMemAccess_CP_742_elements(72) & doMemAccess_CP_742_elements(75);
      gj_doMemAccess_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => doMemAccess_CP_742_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	3 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_sample_completed_
      -- CP-element group 74: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_update_start_
      -- CP-element group 74: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Sample/ack
      -- CP-element group 74: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Update/$entry
      -- CP-element group 74: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Update/req
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_memory_access_lock_822_inst_ack_0, ack => doMemAccess_CP_742_elements(74)); -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => doMemAccess_CP_742_elements(74), ack => WPIPE_memory_access_lock_822_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	82 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	16 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 assign_stmt_640_to_assign_stmt_825/$exit
      -- CP-element group 75: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_update_completed_
      -- CP-element group 75: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Update/$exit
      -- CP-element group 75: 	 assign_stmt_640_to_assign_stmt_825/WPIPE_memory_access_lock_822_Update/ack
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_memory_access_lock_822_inst_ack_1, ack => doMemAccess_CP_742_elements(75)); -- 
    -- CP-element group 76:  place  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	2 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 tag_update_enable
      -- 
    doMemAccess_CP_742_elements(76) <= doMemAccess_CP_742_elements(2);
    -- CP-element group 77:  place  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	3 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 opcode_update_enable
      -- 
    doMemAccess_CP_742_elements(77) <= doMemAccess_CP_742_elements(3);
    -- CP-element group 78:  place  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	4 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 base_addr_update_enable
      -- 
    doMemAccess_CP_742_elements(78) <= doMemAccess_CP_742_elements(4);
    -- CP-element group 79:  place  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	5 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 offset_update_enable
      -- 
    doMemAccess_CP_742_elements(79) <= doMemAccess_CP_742_elements(5);
    -- CP-element group 80:  place  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	6 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 wdata_update_enable
      -- 
    doMemAccess_CP_742_elements(80) <= doMemAccess_CP_742_elements(6);
    -- CP-element group 81:  place  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	7 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 rdata_update_enable
      -- 
    -- CP-element group 82:  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 $exit
      -- 
    doMemAccess_CP_742_elements(82) <= doMemAccess_CP_742_elements(75);
    --  hookup: inputs to control-path 
    doMemAccess_CP_742_elements(81) <= rdata_update_enable;
    -- hookup: output from control-path 
    tag_update_enable <= doMemAccess_CP_742_elements(76);
    opcode_update_enable <= doMemAccess_CP_742_elements(77);
    base_addr_update_enable <= doMemAccess_CP_742_elements(78);
    offset_update_enable <= doMemAccess_CP_742_elements(79);
    wdata_update_enable <= doMemAccess_CP_742_elements(80);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u32_u64_813_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u56_u64_806_wire : std_logic_vector(63 downto 0);
    signal EQ_u3_u1_635_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_638_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_644_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_647_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_653_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_656_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_662_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_665_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_669_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_757_wire : std_logic_vector(0 downto 0);
    signal MUX_732_wire : std_logic_vector(0 downto 0);
    signal MUX_742_742_delayed_1_0_800 : std_logic_vector(63 downto 0);
    signal MUX_744_wire : std_logic_vector(0 downto 0);
    signal MUX_778_wire : std_logic_vector(0 downto 0);
    signal MUX_808_wire : std_logic_vector(63 downto 0);
    signal MUX_815_wire : std_logic_vector(63 downto 0);
    signal OR_u1_u1_666_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_724_724_delayed_17_0_788 : std_logic_vector(0 downto 0);
    signal OR_u64_u64_816_wire : std_logic_vector(63 downto 0);
    signal R_LDB_637_wire_constant : std_logic_vector(2 downto 0);
    signal R_LDD_655_wire_constant : std_logic_vector(2 downto 0);
    signal R_LDSTUB_674_wire_constant : std_logic_vector(2 downto 0);
    signal R_LD_646_wire_constant : std_logic_vector(2 downto 0);
    signal R_LOCKMEM_701_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_696_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_731_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_743_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_777_wire_constant : std_logic_vector(0 downto 0);
    signal R_STB_634_wire_constant : std_logic_vector(2 downto 0);
    signal R_STB_661_wire_constant : std_logic_vector(2 downto 0);
    signal R_STD_652_wire_constant : std_logic_vector(2 downto 0);
    signal R_STD_668_wire_constant : std_logic_vector(2 downto 0);
    signal R_ST_643_wire_constant : std_logic_vector(2 downto 0);
    signal R_ST_664_wire_constant : std_logic_vector(2 downto 0);
    signal R_UNLOCKMEM_702_wire_constant : std_logic_vector(0 downto 0);
    signal R_UNLOCKMEM_728_wire_constant : std_logic_vector(0 downto 0);
    signal R_UNLOCKMEM_740_wire_constant : std_logic_vector(0 downto 0);
    signal R_UNLOCKMEM_774_wire_constant : std_logic_vector(0 downto 0);
    signal R_WRITEMEM_695_wire_constant : std_logic_vector(0 downto 0);
    signal R_WRITEMEM_730_wire_constant : std_logic_vector(0 downto 0);
    signal R_WRITEMEM_742_wire_constant : std_logic_vector(0 downto 0);
    signal R_WRITEMEM_776_wire_constant : std_logic_vector(0 downto 0);
    signal base_addr_716_delayed_17_0_768 : std_logic_vector(63 downto 0);
    signal do_first_byte_692 : std_logic_vector(0 downto 0);
    signal do_ldstub_write_759 : std_logic_vector(0 downto 0);
    signal first_byte_lock_704 : std_logic_vector(0 downto 0);
    signal first_byte_rwbar_698 : std_logic_vector(0 downto 0);
    signal is_byte_access_640 : std_logic_vector(0 downto 0);
    signal is_dword_access_658 : std_logic_vector(0 downto 0);
    signal is_dword_access_739_delayed_16_0_794 : std_logic_vector(0 downto 0);
    signal is_ldstub_664_delayed_1_0_711 : std_logic_vector(0 downto 0);
    signal is_ldstub_676 : std_logic_vector(0 downto 0);
    signal is_ldstub_703_delayed_17_0_752 : std_logic_vector(0 downto 0);
    signal is_ldstub_709_delayed_17_0_762 : std_logic_vector(0 downto 0);
    signal is_word_access_649 : std_logic_vector(0 downto 0);
    signal is_word_access_731_delayed_17_0_791 : std_logic_vector(0 downto 0);
    signal is_write_671 : std_logic_vector(0 downto 0);
    signal konst_756_wire_constant : std_logic_vector(7 downto 0);
    signal konst_781_wire_constant : std_logic_vector(7 downto 0);
    signal konst_798_wire_constant : std_logic_vector(63 downto 0);
    signal konst_807_wire_constant : std_logic_vector(63 downto 0);
    signal konst_814_wire_constant : std_logic_vector(63 downto 0);
    signal mem_lock_707 : std_logic_vector(0 downto 0);
    signal offset_717_delayed_17_0_771 : std_logic_vector(63 downto 0);
    signal r_byte_725 : std_logic_vector(7 downto 0);
    signal r_byte_second_ldstub_783 : std_logic_vector(7 downto 0);
    signal r_dword_749 : std_logic_vector(63 downto 0);
    signal r_word_737 : std_logic_vector(31 downto 0);
    signal tag_710_delayed_17_0_765 : std_logic_vector(7 downto 0);
    signal type_cast_804_wire_constant : std_logic_vector(55 downto 0);
    signal type_cast_811_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(0 downto 0);
    signal w_byte_680 : std_logic_vector(7 downto 0);
    signal w_dword_687 : std_logic_vector(63 downto 0);
    signal w_word_684 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_LDB_637_wire_constant <= "110";
    R_LDD_655_wire_constant <= "101";
    R_LDSTUB_674_wire_constant <= "111";
    R_LD_646_wire_constant <= "100";
    R_LOCKMEM_701_wire_constant <= "1";
    R_READMEM_696_wire_constant <= "1";
    R_READMEM_731_wire_constant <= "1";
    R_READMEM_743_wire_constant <= "1";
    R_READMEM_777_wire_constant <= "1";
    R_STB_634_wire_constant <= "011";
    R_STB_661_wire_constant <= "011";
    R_STD_652_wire_constant <= "010";
    R_STD_668_wire_constant <= "010";
    R_ST_643_wire_constant <= "001";
    R_ST_664_wire_constant <= "001";
    R_UNLOCKMEM_702_wire_constant <= "0";
    R_UNLOCKMEM_728_wire_constant <= "0";
    R_UNLOCKMEM_740_wire_constant <= "0";
    R_UNLOCKMEM_774_wire_constant <= "0";
    R_WRITEMEM_695_wire_constant <= "0";
    R_WRITEMEM_730_wire_constant <= "0";
    R_WRITEMEM_742_wire_constant <= "0";
    R_WRITEMEM_776_wire_constant <= "0";
    konst_756_wire_constant <= "00000000";
    konst_781_wire_constant <= "11111111";
    konst_798_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_807_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_804_wire_constant <= "00000000000000000000000000000000000000000000000000000000";
    type_cast_811_wire_constant <= "00000000000000000000000000000000";
    type_cast_824_wire_constant <= "1";
    -- flow-through select operator MUX_697_inst
    first_byte_rwbar_698 <= R_WRITEMEM_695_wire_constant when (is_write_671(0) /=  '0') else R_READMEM_696_wire_constant;
    -- flow-through select operator MUX_703_inst
    first_byte_lock_704 <= R_LOCKMEM_701_wire_constant when (is_ldstub_676(0) /=  '0') else R_UNLOCKMEM_702_wire_constant;
    -- flow-through select operator MUX_732_inst
    MUX_732_wire <= R_WRITEMEM_730_wire_constant when (is_write_671(0) /=  '0') else R_READMEM_731_wire_constant;
    -- flow-through select operator MUX_744_inst
    MUX_744_wire <= R_WRITEMEM_742_wire_constant when (is_write_671(0) /=  '0') else R_READMEM_743_wire_constant;
    -- flow-through select operator MUX_778_inst
    MUX_778_wire <= R_WRITEMEM_776_wire_constant when (do_ldstub_write_759(0) /=  '0') else R_READMEM_777_wire_constant;
    MUX_799_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_799_inst_req_0;
      MUX_799_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_799_inst_req_1;
      MUX_799_inst_ack_1<= update_ack(0);
      MUX_799_inst: SelectSplitProtocol generic map(name => "MUX_799_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => r_dword_749, y => konst_798_wire_constant, sel => is_dword_access_739_delayed_16_0_794, z => MUX_742_742_delayed_1_0_800, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_808_inst
    MUX_808_wire <= CONCAT_u56_u64_806_wire when (OR_u1_u1_724_724_delayed_17_0_788(0) /=  '0') else konst_807_wire_constant;
    -- flow-through select operator MUX_815_inst
    MUX_815_wire <= CONCAT_u32_u64_813_wire when (is_word_access_731_delayed_17_0_791(0) /=  '0') else konst_814_wire_constant;
    -- flow-through slice operator slice_679_inst
    w_byte_680 <= wdata_buffer(7 downto 0);
    -- flow-through slice operator slice_683_inst
    w_word_684 <= wdata_buffer(31 downto 0);
    W_base_addr_716_delayed_17_0_766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_base_addr_716_delayed_17_0_766_inst_req_0;
      W_base_addr_716_delayed_17_0_766_inst_ack_0<= wack(0);
      rreq(0) <= W_base_addr_716_delayed_17_0_766_inst_req_1;
      W_base_addr_716_delayed_17_0_766_inst_ack_1<= rack(0);
      W_base_addr_716_delayed_17_0_766_inst : InterlockBuffer generic map ( -- 
        name => "W_base_addr_716_delayed_17_0_766_inst",
        buffer_size => 17,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => base_addr_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => base_addr_716_delayed_17_0_768,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_is_dword_access_739_delayed_16_0_792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_is_dword_access_739_delayed_16_0_792_inst_req_0;
      W_is_dword_access_739_delayed_16_0_792_inst_ack_0<= wack(0);
      rreq(0) <= W_is_dword_access_739_delayed_16_0_792_inst_req_1;
      W_is_dword_access_739_delayed_16_0_792_inst_ack_1<= rack(0);
      W_is_dword_access_739_delayed_16_0_792_inst : InterlockBuffer generic map ( -- 
        name => "W_is_dword_access_739_delayed_16_0_792_inst",
        buffer_size => 16,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => is_dword_access_658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => is_dword_access_739_delayed_16_0_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_is_ldstub_664_delayed_1_0_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_is_ldstub_664_delayed_1_0_709_inst_req_0;
      W_is_ldstub_664_delayed_1_0_709_inst_ack_0<= wack(0);
      rreq(0) <= W_is_ldstub_664_delayed_1_0_709_inst_req_1;
      W_is_ldstub_664_delayed_1_0_709_inst_ack_1<= rack(0);
      W_is_ldstub_664_delayed_1_0_709_inst : InterlockBuffer generic map ( -- 
        name => "W_is_ldstub_664_delayed_1_0_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => is_ldstub_676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => is_ldstub_664_delayed_1_0_711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_is_ldstub_703_delayed_17_0_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_is_ldstub_703_delayed_17_0_750_inst_req_0;
      W_is_ldstub_703_delayed_17_0_750_inst_ack_0<= wack(0);
      rreq(0) <= W_is_ldstub_703_delayed_17_0_750_inst_req_1;
      W_is_ldstub_703_delayed_17_0_750_inst_ack_1<= rack(0);
      W_is_ldstub_703_delayed_17_0_750_inst : InterlockBuffer generic map ( -- 
        name => "W_is_ldstub_703_delayed_17_0_750_inst",
        buffer_size => 17,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => is_ldstub_676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => is_ldstub_703_delayed_17_0_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_is_ldstub_709_delayed_17_0_760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_is_ldstub_709_delayed_17_0_760_inst_req_0;
      W_is_ldstub_709_delayed_17_0_760_inst_ack_0<= wack(0);
      rreq(0) <= W_is_ldstub_709_delayed_17_0_760_inst_req_1;
      W_is_ldstub_709_delayed_17_0_760_inst_ack_1<= rack(0);
      W_is_ldstub_709_delayed_17_0_760_inst : InterlockBuffer generic map ( -- 
        name => "W_is_ldstub_709_delayed_17_0_760_inst",
        buffer_size => 17,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => is_ldstub_676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => is_ldstub_709_delayed_17_0_762,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_is_word_access_731_delayed_17_0_789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_is_word_access_731_delayed_17_0_789_inst_req_0;
      W_is_word_access_731_delayed_17_0_789_inst_ack_0<= wack(0);
      rreq(0) <= W_is_word_access_731_delayed_17_0_789_inst_req_1;
      W_is_word_access_731_delayed_17_0_789_inst_ack_1<= rack(0);
      W_is_word_access_731_delayed_17_0_789_inst : InterlockBuffer generic map ( -- 
        name => "W_is_word_access_731_delayed_17_0_789_inst",
        buffer_size => 17,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => is_word_access_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => is_word_access_731_delayed_17_0_791,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_offset_717_delayed_17_0_769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_offset_717_delayed_17_0_769_inst_req_0;
      W_offset_717_delayed_17_0_769_inst_ack_0<= wack(0);
      rreq(0) <= W_offset_717_delayed_17_0_769_inst_req_1;
      W_offset_717_delayed_17_0_769_inst_ack_1<= rack(0);
      W_offset_717_delayed_17_0_769_inst : InterlockBuffer generic map ( -- 
        name => "W_offset_717_delayed_17_0_769_inst",
        buffer_size => 17,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => offset_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => offset_717_delayed_17_0_771,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_tag_710_delayed_17_0_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_tag_710_delayed_17_0_763_inst_req_0;
      W_tag_710_delayed_17_0_763_inst_ack_0<= wack(0);
      rreq(0) <= W_tag_710_delayed_17_0_763_inst_req_1;
      W_tag_710_delayed_17_0_763_inst_ack_1<= rack(0);
      W_tag_710_delayed_17_0_763_inst : InterlockBuffer generic map ( -- 
        name => "W_tag_710_delayed_17_0_763_inst",
        buffer_size => 17,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_710_delayed_17_0_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_w_dword_685_inst
    process(wdata_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := wdata_buffer(63 downto 0);
      w_dword_687 <= tmp_var; -- 
    end process;
    -- flow through binary operator AND_u1_u1_758_inst
    do_ldstub_write_759 <= (is_ldstub_703_delayed_17_0_752 and EQ_u8_u1_757_wire);
    -- flow through binary operator CONCAT_u32_u64_813_inst
    process(type_cast_811_wire_constant, r_word_737) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_811_wire_constant, r_word_737, tmp_var);
      CONCAT_u32_u64_813_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u56_u64_806_inst
    process(type_cast_804_wire_constant, r_byte_725) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_804_wire_constant, r_byte_725, tmp_var);
      CONCAT_u56_u64_806_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_635_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_STB_634_wire_constant, tmp_var);
      EQ_u3_u1_635_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_638_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_LDB_637_wire_constant, tmp_var);
      EQ_u3_u1_638_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_644_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_ST_643_wire_constant, tmp_var);
      EQ_u3_u1_644_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_647_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_LD_646_wire_constant, tmp_var);
      EQ_u3_u1_647_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_653_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_STD_652_wire_constant, tmp_var);
      EQ_u3_u1_653_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_656_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_LDD_655_wire_constant, tmp_var);
      EQ_u3_u1_656_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_662_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_STB_661_wire_constant, tmp_var);
      EQ_u3_u1_662_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_665_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_ST_664_wire_constant, tmp_var);
      EQ_u3_u1_665_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_669_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_STD_668_wire_constant, tmp_var);
      EQ_u3_u1_669_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u3_u1_675_inst
    process(opcode_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(opcode_buffer, R_LDSTUB_674_wire_constant, tmp_var);
      is_ldstub_676 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_757_inst
    process(r_byte_725) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(r_byte_725, konst_756_wire_constant, tmp_var);
      EQ_u8_u1_757_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_639_inst
    is_byte_access_640 <= (EQ_u3_u1_635_wire or EQ_u3_u1_638_wire);
    -- flow through binary operator OR_u1_u1_648_inst
    is_word_access_649 <= (EQ_u3_u1_644_wire or EQ_u3_u1_647_wire);
    -- flow through binary operator OR_u1_u1_657_inst
    is_dword_access_658 <= (EQ_u3_u1_653_wire or EQ_u3_u1_656_wire);
    -- flow through binary operator OR_u1_u1_666_inst
    OR_u1_u1_666_wire <= (EQ_u3_u1_662_wire or EQ_u3_u1_665_wire);
    -- flow through binary operator OR_u1_u1_670_inst
    is_write_671 <= (OR_u1_u1_666_wire or EQ_u3_u1_669_wire);
    -- flow through binary operator OR_u1_u1_691_inst
    do_first_byte_692 <= (is_ldstub_676 or is_byte_access_640);
    -- shared split operator group (20) : OR_u1_u1_787_inst 
    ApIntOr_group_20: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 17);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= is_ldstub_676 & is_byte_access_640;
      OR_u1_u1_724_724_delayed_17_0_788 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u1_u1_787_inst_req_0;
      OR_u1_u1_787_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u1_u1_787_inst_req_1;
      OR_u1_u1_787_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_20_gI: SplitGuardInterface generic map(name => "ApIntOr_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 17,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- flow through binary operator OR_u64_u64_816_inst
    OR_u64_u64_816_wire <= (MUX_808_wire or MUX_815_wire);
    -- flow through binary operator OR_u64_u64_818_inst
    rdata_buffer <= (OR_u64_u64_816_wire or MUX_742_742_delayed_1_0_800);
    -- shared inport operator group (0) : RPIPE_memory_access_lock_706_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_memory_access_lock_706_inst_req_0;
      RPIPE_memory_access_lock_706_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_memory_access_lock_706_inst_req_1;
      RPIPE_memory_access_lock_706_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      mem_lock_707 <= data_out(0 downto 0);
      memory_access_lock_read_0_gI: SplitGuardInterface generic map(name => "memory_access_lock_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      memory_access_lock_read_0: InputPortRevised -- 
        generic map ( name => "memory_access_lock_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => memory_access_lock_pipe_read_req(0),
          oack => memory_access_lock_pipe_read_ack(0),
          odata => memory_access_lock_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_memory_access_lock_713_inst WPIPE_memory_access_lock_822_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_memory_access_lock_713_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_memory_access_lock_822_inst_req_0;
      WPIPE_memory_access_lock_713_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_memory_access_lock_822_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_memory_access_lock_713_inst_req_1;
      update_req_unguarded(0) <= WPIPE_memory_access_lock_822_inst_req_1;
      WPIPE_memory_access_lock_713_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_memory_access_lock_822_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= is_ldstub_676(0);
      guard_vector(1)  <=  not is_ldstub_664_delayed_1_0_711(0);
      data_in <= mem_lock_707 & type_cast_824_wire_constant;
      memory_access_lock_write_0_gI: SplitGuardInterface generic map(name => "memory_access_lock_write_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      memory_access_lock_write_0: OutputPortRevised -- 
        generic map ( name => "memory_access_lock", data_width => 1, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => memory_access_lock_pipe_write_req(0),
          oack => memory_access_lock_pipe_write_ack(0),
          odata => memory_access_lock_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_725_call call_stmt_783_call 
    accessMemoryByteBase_call_group_0: Block -- 
      signal data_in: std_logic_vector(291 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 17, 1 => 17);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_725_call_req_0;
      reqL_unguarded(0) <= call_stmt_783_call_req_0;
      call_stmt_725_call_ack_0 <= ackL_unguarded(1);
      call_stmt_783_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_725_call_req_1;
      reqR_unguarded(0) <= call_stmt_783_call_req_1;
      call_stmt_725_call_ack_1 <= ackR_unguarded(1);
      call_stmt_783_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= is_ldstub_709_delayed_17_0_762(0);
      guard_vector(1)  <= do_first_byte_692(0);
      accessMemoryByteBase_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemoryByteBase_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemoryByteBase_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemoryByteBase_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemoryByteBase_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryByteBase_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & first_byte_lock_704 & first_byte_rwbar_698 & base_addr_buffer & offset_buffer & w_byte_680 & tag_710_delayed_17_0_765 & R_UNLOCKMEM_774_wire_constant & MUX_778_wire & base_addr_716_delayed_17_0_768 & offset_717_delayed_17_0_771 & konst_781_wire_constant;
      r_byte_725 <= data_out(15 downto 8);
      r_byte_second_ldstub_783 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 292,
        owidth => 146,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryByteBase_call_reqs(0),
          ackR => accessMemoryByteBase_call_acks(0),
          dataR => accessMemoryByteBase_call_data(145 downto 0),
          tagR => accessMemoryByteBase_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryByteBase_return_acks(0), -- cross-over
          ackL => accessMemoryByteBase_return_reqs(0), -- cross-over
          dataL => accessMemoryByteBase_return_data(7 downto 0),
          tagL => accessMemoryByteBase_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_737_call 
    accessMemoryWordBase_call_group_1: Block -- 
      signal data_in: std_logic_vector(169 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 17);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_737_call_req_0;
      call_stmt_737_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_737_call_req_1;
      call_stmt_737_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= is_word_access_649(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWordBase_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryWordBase_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_UNLOCKMEM_728_wire_constant & MUX_732_wire & base_addr_buffer & offset_buffer & w_word_684;
      r_word_737 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 170,
        owidth => 170,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWordBase_call_reqs(0),
          ackR => accessMemoryWordBase_call_acks(0),
          dataR => accessMemoryWordBase_call_data(169 downto 0),
          tagR => accessMemoryWordBase_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWordBase_return_acks(0), -- cross-over
          ackL => accessMemoryWordBase_return_reqs(0), -- cross-over
          dataL => accessMemoryWordBase_return_data(31 downto 0),
          tagL => accessMemoryWordBase_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_749_call 
    accessMemoryDwordBase_call_group_2: Block -- 
      signal data_in: std_logic_vector(201 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 16);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_749_call_req_0;
      call_stmt_749_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_749_call_req_1;
      call_stmt_749_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= is_dword_access_658(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDwordBase_call_group_2_gI: SplitGuardInterface generic map(name => "accessMemoryDwordBase_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_UNLOCKMEM_740_wire_constant & MUX_744_wire & base_addr_buffer & offset_buffer & w_dword_687;
      r_dword_749 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 202,
        owidth => 202,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDwordBase_call_reqs(0),
          ackR => accessMemoryDwordBase_call_acks(0),
          dataR => accessMemoryDwordBase_call_data(201 downto 0),
          tagR => accessMemoryDwordBase_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDwordBase_return_acks(0), -- cross-over
          ackL => accessMemoryDwordBase_return_reqs(0), -- cross-over
          dataL => accessMemoryDwordBase_return_data(63 downto 0),
          tagL => accessMemoryDwordBase_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end doMemAccess_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getBaseIndex_Volatile is -- 
  port ( -- 
    queue_type : in  std_logic_vector(1 downto 0);
    server_id : in  std_logic_vector(7 downto 0);
    base_index : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity getBaseIndex_Volatile;
architecture getBaseIndex_Volatile_arch of getBaseIndex_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(10-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal queue_type_buffer :  std_logic_vector(1 downto 0);
  signal server_id_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal base_index_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  queue_type_buffer <= queue_type;
  server_id_buffer <= server_id;
  -- output handling  -------------------------------------------------------
  base_index <= base_index_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_141_wire : std_logic_vector(7 downto 0);
    signal ADD_u8_u8_152_wire : std_logic_vector(7 downto 0);
    signal EQ_u2_u1_130_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_136_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_147_wire : std_logic_vector(0 downto 0);
    signal MUL_u8_u8_140_wire : std_logic_vector(7 downto 0);
    signal MUL_u8_u8_151_wire : std_logic_vector(7 downto 0);
    signal MUX_133_wire : std_logic_vector(7 downto 0);
    signal MUX_143_wire : std_logic_vector(7 downto 0);
    signal MUX_154_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_144_wire : std_logic_vector(7 downto 0);
    signal R_FREEQUEUE_129_wire_constant : std_logic_vector(1 downto 0);
    signal R_RXQUEUE_146_wire_constant : std_logic_vector(1 downto 0);
    signal R_TXQUEUE_135_wire_constant : std_logic_vector(1 downto 0);
    signal konst_131_wire_constant : std_logic_vector(7 downto 0);
    signal konst_132_wire_constant : std_logic_vector(7 downto 0);
    signal konst_137_wire_constant : std_logic_vector(7 downto 0);
    signal konst_139_wire_constant : std_logic_vector(7 downto 0);
    signal konst_142_wire_constant : std_logic_vector(7 downto 0);
    signal konst_148_wire_constant : std_logic_vector(7 downto 0);
    signal konst_150_wire_constant : std_logic_vector(7 downto 0);
    signal konst_153_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_FREEQUEUE_129_wire_constant <= "00";
    R_RXQUEUE_146_wire_constant <= "10";
    R_TXQUEUE_135_wire_constant <= "01";
    konst_131_wire_constant <= "11001000";
    konst_132_wire_constant <= "00000000";
    konst_137_wire_constant <= "10000000";
    konst_139_wire_constant <= "00001000";
    konst_142_wire_constant <= "00000000";
    konst_148_wire_constant <= "00001000";
    konst_150_wire_constant <= "00001000";
    konst_153_wire_constant <= "00000000";
    -- flow-through select operator MUX_133_inst
    MUX_133_wire <= konst_131_wire_constant when (EQ_u2_u1_130_wire(0) /=  '0') else konst_132_wire_constant;
    -- flow-through select operator MUX_143_inst
    MUX_143_wire <= ADD_u8_u8_141_wire when (EQ_u2_u1_136_wire(0) /=  '0') else konst_142_wire_constant;
    -- flow-through select operator MUX_154_inst
    MUX_154_wire <= ADD_u8_u8_152_wire when (EQ_u2_u1_147_wire(0) /=  '0') else konst_153_wire_constant;
    -- flow through binary operator ADD_u8_u8_141_inst
    ADD_u8_u8_141_wire <= std_logic_vector(unsigned(MUL_u8_u8_140_wire) + unsigned(konst_137_wire_constant));
    -- flow through binary operator ADD_u8_u8_152_inst
    ADD_u8_u8_152_wire <= std_logic_vector(unsigned(MUL_u8_u8_151_wire) + unsigned(konst_148_wire_constant));
    -- flow through binary operator EQ_u2_u1_130_inst
    process(queue_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(queue_type_buffer, R_FREEQUEUE_129_wire_constant, tmp_var);
      EQ_u2_u1_130_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_136_inst
    process(queue_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(queue_type_buffer, R_TXQUEUE_135_wire_constant, tmp_var);
      EQ_u2_u1_136_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_147_inst
    process(queue_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(queue_type_buffer, R_RXQUEUE_146_wire_constant, tmp_var);
      EQ_u2_u1_147_wire <= tmp_var; --
    end process;
    -- flow through binary operator MUL_u8_u8_140_inst
    process(server_id_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(server_id_buffer, konst_139_wire_constant, tmp_var);
      MUL_u8_u8_140_wire <= tmp_var; --
    end process;
    -- flow through binary operator MUL_u8_u8_151_inst
    process(server_id_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(server_id_buffer, konst_150_wire_constant, tmp_var);
      MUL_u8_u8_151_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u8_u8_144_inst
    OR_u8_u8_144_wire <= (MUX_133_wire or MUX_143_wire);
    -- flow through binary operator OR_u8_u8_155_inst
    base_index_buffer <= (OR_u8_u8_144_wire or MUX_154_wire);
    -- 
  end Block; -- data_path
  -- 
end getBaseIndex_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getQueueBufPointer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_type : in  std_logic_vector(1 downto 0);
    server_id : in  std_logic_vector(7 downto 0);
    qptr : out  std_logic_vector(63 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_call_acks : in   std_logic_vector(0 downto 0);
    accessRegister_call_data : out  std_logic_vector(44 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_return_acks : in   std_logic_vector(0 downto 0);
    accessRegister_return_data : in   std_logic_vector(31 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueBufPointer;
architecture getQueueBufPointer_arch of getQueueBufPointer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 10)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_type_buffer :  std_logic_vector(1 downto 0);
  signal queue_type_update_enable: Boolean;
  signal server_id_buffer :  std_logic_vector(7 downto 0);
  signal server_id_update_enable: Boolean;
  -- output port buffer signals
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal getQueueBufPointer_CP_1416_start: Boolean;
  signal getQueueBufPointer_CP_1416_symbol: Boolean;
  -- volatile/operator module components. 
  component getBaseIndex_Volatile is -- 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      base_index : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1057_call_ack_0 : boolean;
  signal call_stmt_1057_call_ack_1 : boolean;
  signal W_base_idx_1044_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1070_inst_req_0 : boolean;
  signal call_stmt_1057_call_req_0 : boolean;
  signal CONCAT_u32_u64_1070_inst_ack_0 : boolean;
  signal call_stmt_1057_call_req_1 : boolean;
  signal CONCAT_u32_u64_1070_inst_ack_1 : boolean;
  signal W_base_idx_1044_inst_ack_0 : boolean;
  signal W_base_idx_1044_inst_req_1 : boolean;
  signal W_base_idx_1044_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1070_inst_req_1 : boolean;
  signal call_stmt_1066_call_ack_1 : boolean;
  signal call_stmt_1066_call_req_1 : boolean;
  signal call_stmt_1066_call_ack_0 : boolean;
  signal call_stmt_1066_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueBufPointer_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 10) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(1 downto 0) <= queue_type;
  queue_type_buffer <= in_buffer_data_out(1 downto 0);
  in_buffer_data_in(9 downto 2) <= server_id;
  server_id_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(tag_length + 9 downto 10) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 9 downto 10);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueBufPointer_CP_1416_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueBufPointer_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= qptr_buffer;
  qptr <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueBufPointer_CP_1416_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueBufPointer_CP_1416_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueBufPointer_CP_1416_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueBufPointer_CP_1416: Block -- control-path 
    signal getQueueBufPointer_CP_1416_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    getQueueBufPointer_CP_1416_elements(0) <= getQueueBufPointer_CP_1416_start;
    getQueueBufPointer_CP_1416_symbol <= getQueueBufPointer_CP_1416_elements(10);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_update_start_
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_update_start_
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Sample/req
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_sample_start_
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Update/req
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_update_start_
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Update/cr
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/$entry
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_update_start_
      -- CP-element group 0: 	 $entry
      -- 
    req_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(0), ack => W_base_idx_1044_inst_req_0); -- 
    req_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(0), ack => W_base_idx_1044_inst_req_1); -- 
    ccr_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(0), ack => call_stmt_1057_call_req_1); -- 
    ccr_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(0), ack => call_stmt_1066_call_req_1); -- 
    cr_1476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(0), ack => CONCAT_u32_u64_1070_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Sample/ack
      -- 
    ack_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_idx_1044_inst_ack_0, ack => getQueueBufPointer_CP_1416_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Sample/crr
      -- CP-element group 2: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_update_completed_
      -- CP-element group 2: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1048_to_assign_stmt_1071/assign_stmt_1048_Update/ack
      -- CP-element group 2: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_sample_start_
      -- CP-element group 2: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Sample/$entry
      -- 
    ack_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_idx_1044_inst_ack_1, ack => getQueueBufPointer_CP_1416_elements(2)); -- 
    crr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(2), ack => call_stmt_1057_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Sample/cra
      -- CP-element group 3: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_sample_completed_
      -- 
    cra_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1057_call_ack_0, ack => getQueueBufPointer_CP_1416_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Update/cca
      -- CP-element group 4: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_Update/$exit
      -- CP-element group 4: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_update_completed_
      -- 
    cca_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1057_call_ack_1, ack => getQueueBufPointer_CP_1416_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_sample_start_
      -- CP-element group 5: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Sample/crr
      -- CP-element group 5: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Sample/$entry
      -- 
    crr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(5), ack => call_stmt_1066_call_req_0); -- 
    getQueueBufPointer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "getQueueBufPointer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getQueueBufPointer_CP_1416_elements(2) & getQueueBufPointer_CP_1416_elements(11);
      gj_getQueueBufPointer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getQueueBufPointer_CP_1416_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_sample_completed_
      -- CP-element group 6: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Sample/cra
      -- CP-element group 6: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Sample/$exit
      -- 
    cra_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1066_call_ack_0, ack => getQueueBufPointer_CP_1416_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_update_completed_
      -- CP-element group 7: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Update/cca
      -- CP-element group 7: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1066_Update/$exit
      -- 
    cca_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1066_call_ack_1, ack => getQueueBufPointer_CP_1416_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Sample/rr
      -- CP-element group 8: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_sample_start_
      -- 
    rr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueBufPointer_CP_1416_elements(8), ack => CONCAT_u32_u64_1070_inst_req_0); -- 
    getQueueBufPointer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "getQueueBufPointer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getQueueBufPointer_CP_1416_elements(4) & getQueueBufPointer_CP_1416_elements(7);
      gj_getQueueBufPointer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getQueueBufPointer_CP_1416_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_sample_completed_
      -- CP-element group 9: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Sample/ra
      -- 
    ra_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1070_inst_ack_0, ack => getQueueBufPointer_CP_1416_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_update_completed_
      -- CP-element group 10: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Update/ca
      -- CP-element group 10: 	 assign_stmt_1048_to_assign_stmt_1071/$exit
      -- CP-element group 10: 	 assign_stmt_1048_to_assign_stmt_1071/CONCAT_u32_u64_1070_Update/$exit
      -- CP-element group 10: 	 $exit
      -- 
    ca_1477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1070_inst_ack_1, ack => getQueueBufPointer_CP_1416_elements(10)); -- 
    -- CP-element group 11:  transition  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	4 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 assign_stmt_1048_to_assign_stmt_1071/call_stmt_1057_call_stmt_1066_delay
      -- 
    -- Element group getQueueBufPointer_CP_1416_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => getQueueBufPointer_CP_1416_elements(4), ack => getQueueBufPointer_CP_1416_elements(11), clk => clk, reset =>reset);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_1053_wire : std_logic_vector(7 downto 0);
    signal ADD_u8_u8_1062_wire : std_logic_vector(7 downto 0);
    signal R_READMEM_1049_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_1058_wire_constant : std_logic_vector(0 downto 0);
    signal base_idx_1048 : std_logic_vector(7 downto 0);
    signal call_getBaseIndex_expr_1047_wire : std_logic_vector(7 downto 0);
    signal konst_1050_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1052_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1059_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1061_wire_constant : std_logic_vector(7 downto 0);
    signal qptr_h_1057 : std_logic_vector(31 downto 0);
    signal qptr_l_1066 : std_logic_vector(31 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_1049_wire_constant <= "1";
    R_READMEM_1058_wire_constant <= "1";
    konst_1050_wire_constant <= "1111";
    konst_1052_wire_constant <= "00000100";
    konst_1059_wire_constant <= "1111";
    konst_1061_wire_constant <= "00000101";
    type_cast_1055_wire_constant <= "00000000000000000000000000000000";
    type_cast_1064_wire_constant <= "00000000000000000000000000000000";
    W_base_idx_1044_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_base_idx_1044_inst_req_0;
      W_base_idx_1044_inst_ack_0<= wack(0);
      rreq(0) <= W_base_idx_1044_inst_req_1;
      W_base_idx_1044_inst_ack_1<= rack(0);
      W_base_idx_1044_inst : InterlockBuffer generic map ( -- 
        name => "W_base_idx_1044_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_getBaseIndex_expr_1047_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => base_idx_1048,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- flow through binary operator ADD_u8_u8_1053_inst
    ADD_u8_u8_1053_wire <= std_logic_vector(unsigned(base_idx_1048) + unsigned(konst_1052_wire_constant));
    -- flow through binary operator ADD_u8_u8_1062_inst
    ADD_u8_u8_1062_wire <= std_logic_vector(unsigned(base_idx_1048) + unsigned(konst_1061_wire_constant));
    -- shared split operator group (2) : CONCAT_u32_u64_1070_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= qptr_h_1057 & qptr_l_1066;
      qptr_buffer <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1070_inst_req_0;
      CONCAT_u32_u64_1070_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1070_inst_req_1;
      CONCAT_u32_u64_1070_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    volatile_operator_getBaseIndex_2364: getBaseIndex_Volatile port map(queue_type => queue_type_buffer, server_id => server_id_buffer, base_index => call_getBaseIndex_expr_1047_wire); 
    -- shared call operator group (1) : call_stmt_1066_call call_stmt_1057_call 
    accessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1066_call_req_0;
      reqL_unguarded(0) <= call_stmt_1057_call_req_0;
      call_stmt_1066_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1057_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1066_call_req_1;
      reqR_unguarded(0) <= call_stmt_1057_call_req_1;
      call_stmt_1066_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1057_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessRegister_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "accessRegister_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "accessRegister_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_READMEM_1058_wire_constant & konst_1059_wire_constant & ADD_u8_u8_1062_wire & type_cast_1064_wire_constant & R_READMEM_1049_wire_constant & konst_1050_wire_constant & ADD_u8_u8_1053_wire & type_cast_1055_wire_constant;
      qptr_l_1066 <= data_out(63 downto 32);
      qptr_h_1057 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 90,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getQueueBufPointer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    buf_base_addr : in  std_logic_vector(63 downto 0);
    read_index : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(63 downto 0);
    accessQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueElement_call_data : out  std_logic_vector(168 downto 0);
    accessQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueElement_return_data : in   std_logic_vector(63 downto 0);
    accessQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal buf_base_addr_buffer :  std_logic_vector(63 downto 0);
  signal buf_base_addr_update_enable: Boolean;
  signal read_index_buffer :  std_logic_vector(31 downto 0);
  signal read_index_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(63 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_1537_start: Boolean;
  signal getQueueElement_CP_1537_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      index : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1128_call_req_1 : boolean;
  signal call_stmt_1128_call_ack_1 : boolean;
  signal call_stmt_1128_call_ack_0 : boolean;
  signal call_stmt_1128_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= buf_base_addr;
  buf_base_addr_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(103 downto 72) <= read_index;
  read_index_buffer <= in_buffer_data_out(103 downto 72);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_1537_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_1537_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_1537_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_1537_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_1537: Block -- control-path 
    signal getQueueElement_CP_1537_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_1537_elements(0) <= getQueueElement_CP_1537_start;
    getQueueElement_CP_1537_symbol <= getQueueElement_CP_1537_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_1128/call_stmt_1128_Update/ccr
      -- CP-element group 0: 	 call_stmt_1128/call_stmt_1128_Update/$entry
      -- CP-element group 0: 	 call_stmt_1128/call_stmt_1128_Sample/crr
      -- CP-element group 0: 	 call_stmt_1128/call_stmt_1128_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1128/call_stmt_1128_update_start_
      -- CP-element group 0: 	 call_stmt_1128/call_stmt_1128_sample_start_
      -- CP-element group 0: 	 call_stmt_1128/$entry
      -- CP-element group 0: 	 $entry
      -- 
    ccr_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_1537_elements(0), ack => call_stmt_1128_call_req_1); -- 
    crr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_1537_elements(0), ack => call_stmt_1128_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1128/call_stmt_1128_Sample/cra
      -- CP-element group 1: 	 call_stmt_1128/call_stmt_1128_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1128/call_stmt_1128_sample_completed_
      -- 
    cra_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1128_call_ack_0, ack => getQueueElement_CP_1537_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_1128/call_stmt_1128_Update/cca
      -- CP-element group 2: 	 call_stmt_1128/call_stmt_1128_Update/$exit
      -- CP-element group 2: 	 call_stmt_1128/call_stmt_1128_update_completed_
      -- CP-element group 2: 	 call_stmt_1128/$exit
      -- CP-element group 2: 	 $exit
      -- 
    cca_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1128_call_ack_1, ack => getQueueElement_CP_1537_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_READMEM_1122_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1126_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    R_READMEM_1122_wire_constant <= "1";
    type_cast_1126_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_1128_call 
    accessQueueElement_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1128_call_req_0;
      call_stmt_1128_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1128_call_req_1;
      call_stmt_1128_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueElement_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueElement_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_1122_wire_constant & buf_base_addr_buffer & read_index_buffer & type_cast_1126_wire_constant;
      q_r_data_buffer <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueElement_call_reqs(0),
          ackR => accessQueueElement_call_acks(0),
          dataR => accessQueueElement_call_data(168 downto 0),
          tagR => accessQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueElement_return_acks(0), -- cross-over
          ackL => accessQueueElement_return_reqs(0), -- cross-over
          dataL => accessQueueElement_return_data(63 downto 0),
          tagL => accessQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getQueueLength is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    q_base_address : in  std_logic_vector(63 downto 0);
    queue_length : out  std_logic_vector(31 downto 0);
    accessQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueLength_call_data : out  std_logic_vector(104 downto 0);
    accessQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueLength_return_data : in   std_logic_vector(31 downto 0);
    accessQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueLength;
architecture getQueueLength_arch of getQueueLength is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(63 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal queue_length_buffer :  std_logic_vector(31 downto 0);
  signal queue_length_update_enable: Boolean;
  signal getQueueLength_CP_1356_start: Boolean;
  signal getQueueLength_CP_1356_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1012_call_req_0 : boolean;
  signal call_stmt_1012_call_ack_0 : boolean;
  signal call_stmt_1012_call_req_1 : boolean;
  signal call_stmt_1012_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueLength_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueLength_CP_1356_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueLength_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= queue_length_buffer;
  queue_length <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_1356_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueLength_CP_1356_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_1356_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueLength_CP_1356: Block -- control-path 
    signal getQueueLength_CP_1356_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    getQueueLength_CP_1356_elements(0) <= getQueueLength_CP_1356_start;
    getQueueLength_CP_1356_symbol <= getQueueLength_CP_1356_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1012/$entry
      -- CP-element group 0: 	 call_stmt_1012/call_stmt_1012_sample_start_
      -- CP-element group 0: 	 call_stmt_1012/call_stmt_1012_update_start_
      -- CP-element group 0: 	 call_stmt_1012/call_stmt_1012_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1012/call_stmt_1012_Sample/crr
      -- CP-element group 0: 	 call_stmt_1012/call_stmt_1012_Update/$entry
      -- CP-element group 0: 	 call_stmt_1012/call_stmt_1012_Update/ccr
      -- 
    crr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_1356_elements(0), ack => call_stmt_1012_call_req_0); -- 
    ccr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_1356_elements(0), ack => call_stmt_1012_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1012/call_stmt_1012_sample_completed_
      -- CP-element group 1: 	 call_stmt_1012/call_stmt_1012_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1012/call_stmt_1012_Sample/cra
      -- 
    cra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1012_call_ack_0, ack => getQueueLength_CP_1356_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1012/$exit
      -- CP-element group 2: 	 call_stmt_1012/call_stmt_1012_update_completed_
      -- CP-element group 2: 	 call_stmt_1012/call_stmt_1012_Update/$exit
      -- CP-element group 2: 	 call_stmt_1012/call_stmt_1012_Update/cca
      -- 
    cca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1012_call_ack_1, ack => getQueueLength_CP_1356_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_READMEM_1007_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_1007_wire_constant <= "1";
    type_cast_1010_wire_constant <= "00000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_1012_call 
    accessQueueLength_call_group_0: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1012_call_req_0;
      call_stmt_1012_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1012_call_req_1;
      call_stmt_1012_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueLength_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueLength_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_1007_wire_constant & q_base_address_buffer & type_cast_1010_wire_constant;
      queue_length_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueLength_call_reqs(0),
          ackR => accessQueueLength_call_acks(0),
          dataR => accessQueueLength_call_data(104 downto 0),
          tagR => accessQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueLength_return_acks(0), -- cross-over
          ackL => accessQueueLength_return_reqs(0), -- cross-over
          dataL => accessQueueLength_return_data(31 downto 0),
          tagL => accessQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueLength_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getQueueLockPointer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_type : in  std_logic_vector(1 downto 0);
    server_id : in  std_logic_vector(7 downto 0);
    qptr : out  std_logic_vector(63 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_call_acks : in   std_logic_vector(0 downto 0);
    accessRegister_call_data : out  std_logic_vector(44 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_return_acks : in   std_logic_vector(0 downto 0);
    accessRegister_return_data : in   std_logic_vector(31 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueLockPointer;
architecture getQueueLockPointer_arch of getQueueLockPointer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 10)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_type_buffer :  std_logic_vector(1 downto 0);
  signal queue_type_update_enable: Boolean;
  signal server_id_buffer :  std_logic_vector(7 downto 0);
  signal server_id_update_enable: Boolean;
  -- output port buffer signals
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal getQueueLockPointer_CP_1079_start: Boolean;
  signal getQueueLockPointer_CP_1079_symbol: Boolean;
  -- volatile/operator module components. 
  component getBaseIndex_Volatile is -- 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      base_index : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_892_call_ack_1 : boolean;
  signal call_stmt_883_call_req_0 : boolean;
  signal CONCAT_u32_u64_896_inst_req_0 : boolean;
  signal call_stmt_892_call_req_1 : boolean;
  signal call_stmt_883_call_req_1 : boolean;
  signal call_stmt_883_call_ack_0 : boolean;
  signal CONCAT_u32_u64_896_inst_ack_0 : boolean;
  signal call_stmt_892_call_req_0 : boolean;
  signal CONCAT_u32_u64_896_inst_ack_1 : boolean;
  signal call_stmt_883_call_ack_1 : boolean;
  signal CONCAT_u32_u64_896_inst_req_1 : boolean;
  signal W_base_idx_870_inst_ack_1 : boolean;
  signal W_base_idx_870_inst_req_1 : boolean;
  signal W_base_idx_870_inst_ack_0 : boolean;
  signal W_base_idx_870_inst_req_0 : boolean;
  signal call_stmt_892_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueLockPointer_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 10) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(1 downto 0) <= queue_type;
  queue_type_buffer <= in_buffer_data_out(1 downto 0);
  in_buffer_data_in(9 downto 2) <= server_id;
  server_id_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(tag_length + 9 downto 10) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 9 downto 10);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueLockPointer_CP_1079_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueLockPointer_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= qptr_buffer;
  qptr <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLockPointer_CP_1079_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueLockPointer_CP_1079_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLockPointer_CP_1079_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueLockPointer_CP_1079: Block -- control-path 
    signal getQueueLockPointer_CP_1079_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    getQueueLockPointer_CP_1079_elements(0) <= getQueueLockPointer_CP_1079_start;
    getQueueLockPointer_CP_1079_symbol <= getQueueLockPointer_CP_1079_elements(10);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Update/ccr
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/$entry
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Update/ccr
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_update_start_
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Update/$entry
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Update/$entry
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_update_start_
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_sample_start_
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_update_start_
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Update/cr
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Update/req
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Update/$entry
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Sample/req
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_update_start_
      -- 
    req_1092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(0), ack => W_base_idx_870_inst_req_0); -- 
    req_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(0), ack => W_base_idx_870_inst_req_1); -- 
    ccr_1111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(0), ack => call_stmt_883_call_req_1); -- 
    ccr_1125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(0), ack => call_stmt_892_call_req_1); -- 
    cr_1139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(0), ack => CONCAT_u32_u64_896_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_sample_completed_
      -- CP-element group 1: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Sample/ack
      -- CP-element group 1: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Sample/$exit
      -- 
    ack_1093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_idx_870_inst_ack_0, ack => getQueueLockPointer_CP_1079_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Sample/crr
      -- CP-element group 2: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_sample_start_
      -- CP-element group 2: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Update/ack
      -- CP-element group 2: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_Update/$exit
      -- CP-element group 2: 	 assign_stmt_874_to_assign_stmt_897/assign_stmt_874_update_completed_
      -- 
    ack_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_idx_870_inst_ack_1, ack => getQueueLockPointer_CP_1079_elements(2)); -- 
    crr_1106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(2), ack => call_stmt_883_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Sample/cra
      -- CP-element group 3: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_sample_completed_
      -- 
    cra_1107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_883_call_ack_0, ack => getQueueLockPointer_CP_1079_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Update/$exit
      -- CP-element group 4: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_update_completed_
      -- CP-element group 4: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_Update/cca
      -- 
    cca_1112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_883_call_ack_1, ack => getQueueLockPointer_CP_1079_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_sample_start_
      -- CP-element group 5: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Sample/crr
      -- 
    crr_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(5), ack => call_stmt_892_call_req_0); -- 
    getQueueLockPointer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "getQueueLockPointer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getQueueLockPointer_CP_1079_elements(2) & getQueueLockPointer_CP_1079_elements(11);
      gj_getQueueLockPointer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getQueueLockPointer_CP_1079_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_sample_completed_
      -- CP-element group 6: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Sample/cra
      -- 
    cra_1121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_892_call_ack_0, ack => getQueueLockPointer_CP_1079_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Update/cca
      -- CP-element group 7: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_update_completed_
      -- CP-element group 7: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_892_Update/$exit
      -- 
    cca_1126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_892_call_ack_1, ack => getQueueLockPointer_CP_1079_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Sample/rr
      -- CP-element group 8: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_sample_start_
      -- 
    rr_1134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLockPointer_CP_1079_elements(8), ack => CONCAT_u32_u64_896_inst_req_0); -- 
    getQueueLockPointer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "getQueueLockPointer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getQueueLockPointer_CP_1079_elements(4) & getQueueLockPointer_CP_1079_elements(7);
      gj_getQueueLockPointer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getQueueLockPointer_CP_1079_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Sample/ra
      -- CP-element group 9: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_sample_completed_
      -- 
    ra_1135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_896_inst_ack_0, ack => getQueueLockPointer_CP_1079_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_874_to_assign_stmt_897/$exit
      -- CP-element group 10: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Update/ca
      -- CP-element group 10: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_Update/$exit
      -- CP-element group 10: 	 assign_stmt_874_to_assign_stmt_897/CONCAT_u32_u64_896_update_completed_
      -- CP-element group 10: 	 $exit
      -- 
    ca_1140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_896_inst_ack_1, ack => getQueueLockPointer_CP_1079_elements(10)); -- 
    -- CP-element group 11:  transition  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	4 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 assign_stmt_874_to_assign_stmt_897/call_stmt_883_call_stmt_892_delay
      -- 
    -- Element group getQueueLockPointer_CP_1079_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => getQueueLockPointer_CP_1079_elements(4), ack => getQueueLockPointer_CP_1079_elements(11), clk => clk, reset =>reset);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_879_wire : std_logic_vector(7 downto 0);
    signal ADD_u8_u8_888_wire : std_logic_vector(7 downto 0);
    signal R_READMEM_875_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_884_wire_constant : std_logic_vector(0 downto 0);
    signal base_idx_874 : std_logic_vector(7 downto 0);
    signal call_getBaseIndex_expr_873_wire : std_logic_vector(7 downto 0);
    signal konst_876_wire_constant : std_logic_vector(3 downto 0);
    signal konst_878_wire_constant : std_logic_vector(7 downto 0);
    signal konst_885_wire_constant : std_logic_vector(3 downto 0);
    signal konst_887_wire_constant : std_logic_vector(7 downto 0);
    signal qptr_h_883 : std_logic_vector(31 downto 0);
    signal qptr_l_892 : std_logic_vector(31 downto 0);
    signal type_cast_881_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_875_wire_constant <= "1";
    R_READMEM_884_wire_constant <= "1";
    konst_876_wire_constant <= "1111";
    konst_878_wire_constant <= "00000010";
    konst_885_wire_constant <= "1111";
    konst_887_wire_constant <= "00000011";
    type_cast_881_wire_constant <= "00000000000000000000000000000000";
    type_cast_890_wire_constant <= "00000000000000000000000000000000";
    W_base_idx_870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_base_idx_870_inst_req_0;
      W_base_idx_870_inst_ack_0<= wack(0);
      rreq(0) <= W_base_idx_870_inst_req_1;
      W_base_idx_870_inst_ack_1<= rack(0);
      W_base_idx_870_inst : InterlockBuffer generic map ( -- 
        name => "W_base_idx_870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_getBaseIndex_expr_873_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => base_idx_874,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- flow through binary operator ADD_u8_u8_879_inst
    ADD_u8_u8_879_wire <= std_logic_vector(unsigned(base_idx_874) + unsigned(konst_878_wire_constant));
    -- flow through binary operator ADD_u8_u8_888_inst
    ADD_u8_u8_888_wire <= std_logic_vector(unsigned(base_idx_874) + unsigned(konst_887_wire_constant));
    -- shared split operator group (2) : CONCAT_u32_u64_896_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= qptr_h_883 & qptr_l_892;
      qptr_buffer <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_896_inst_req_0;
      CONCAT_u32_u64_896_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_896_inst_req_1;
      CONCAT_u32_u64_896_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    volatile_operator_getBaseIndex_1889: getBaseIndex_Volatile port map(queue_type => queue_type_buffer, server_id => server_id_buffer, base_index => call_getBaseIndex_expr_873_wire); 
    -- shared call operator group (1) : call_stmt_892_call call_stmt_883_call 
    accessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_892_call_req_0;
      reqL_unguarded(0) <= call_stmt_883_call_req_0;
      call_stmt_892_call_ack_0 <= ackL_unguarded(1);
      call_stmt_883_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_892_call_req_1;
      reqR_unguarded(0) <= call_stmt_883_call_req_1;
      call_stmt_892_call_ack_1 <= ackR_unguarded(1);
      call_stmt_883_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessRegister_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "accessRegister_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "accessRegister_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_READMEM_884_wire_constant & konst_885_wire_constant & ADD_u8_u8_888_wire & type_cast_890_wire_constant & R_READMEM_875_wire_constant & konst_876_wire_constant & ADD_u8_u8_879_wire & type_cast_881_wire_constant;
      qptr_l_892 <= data_out(63 downto 32);
      qptr_h_883 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 90,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getQueueLockPointer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getQueuePointer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_type : in  std_logic_vector(1 downto 0);
    server_id : in  std_logic_vector(7 downto 0);
    qptr : out  std_logic_vector(63 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_call_acks : in   std_logic_vector(0 downto 0);
    accessRegister_call_data : out  std_logic_vector(44 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_return_acks : in   std_logic_vector(0 downto 0);
    accessRegister_return_data : in   std_logic_vector(31 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointer;
architecture getQueuePointer_arch of getQueuePointer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 10)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_type_buffer :  std_logic_vector(1 downto 0);
  signal queue_type_update_enable: Boolean;
  signal server_id_buffer :  std_logic_vector(7 downto 0);
  signal server_id_update_enable: Boolean;
  -- output port buffer signals
  signal qptr_buffer :  std_logic_vector(63 downto 0);
  signal qptr_update_enable: Boolean;
  signal getQueuePointer_CP_134_start: Boolean;
  signal getQueuePointer_CP_134_symbol: Boolean;
  -- volatile/operator module components. 
  component getBaseIndex_Volatile is -- 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      base_index : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_base_idx_247_inst_req_0 : boolean;
  signal W_base_idx_247_inst_ack_0 : boolean;
  signal W_base_idx_247_inst_req_1 : boolean;
  signal W_base_idx_247_inst_ack_1 : boolean;
  signal call_stmt_258_call_req_0 : boolean;
  signal call_stmt_258_call_ack_0 : boolean;
  signal call_stmt_258_call_req_1 : boolean;
  signal call_stmt_258_call_ack_1 : boolean;
  signal call_stmt_267_call_req_0 : boolean;
  signal call_stmt_267_call_ack_0 : boolean;
  signal call_stmt_267_call_req_1 : boolean;
  signal call_stmt_267_call_ack_1 : boolean;
  signal CONCAT_u32_u64_271_inst_req_0 : boolean;
  signal CONCAT_u32_u64_271_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_271_inst_req_1 : boolean;
  signal CONCAT_u32_u64_271_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointer_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 10) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(1 downto 0) <= queue_type;
  queue_type_buffer <= in_buffer_data_out(1 downto 0);
  in_buffer_data_in(9 downto 2) <= server_id;
  server_id_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(tag_length + 9 downto 10) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 9 downto 10);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointer_CP_134_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointer_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= qptr_buffer;
  qptr <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointer_CP_134_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointer_CP_134_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointer_CP_134_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointer_CP_134: Block -- control-path 
    signal getQueuePointer_CP_134_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    getQueuePointer_CP_134_elements(0) <= getQueuePointer_CP_134_start;
    getQueuePointer_CP_134_symbol <= getQueuePointer_CP_134_elements(10);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/$entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_sample_start_
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_update_start_
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Sample/req
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Update/$entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Update/req
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_update_start_
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Update/$entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Update/ccr
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_update_start_
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Update/$entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Update/ccr
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_update_start_
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Update/$entry
      -- CP-element group 0: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Update/cr
      -- 
    req_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(0), ack => W_base_idx_247_inst_req_0); -- 
    req_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(0), ack => W_base_idx_247_inst_req_1); -- 
    ccr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(0), ack => call_stmt_258_call_req_1); -- 
    ccr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(0), ack => call_stmt_267_call_req_1); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(0), ack => CONCAT_u32_u64_271_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_sample_completed_
      -- CP-element group 1: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Sample/ack
      -- 
    ack_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_idx_247_inst_ack_0, ack => getQueuePointer_CP_134_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_update_completed_
      -- CP-element group 2: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Update/$exit
      -- CP-element group 2: 	 assign_stmt_251_to_assign_stmt_272/assign_stmt_251_Update/ack
      -- CP-element group 2: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_sample_start_
      -- CP-element group 2: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Sample/crr
      -- 
    ack_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_base_idx_247_inst_ack_1, ack => getQueuePointer_CP_134_elements(2)); -- 
    crr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(2), ack => call_stmt_258_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_sample_completed_
      -- CP-element group 3: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Sample/cra
      -- 
    cra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_258_call_ack_0, ack => getQueuePointer_CP_134_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_update_completed_
      -- CP-element group 4: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Update/$exit
      -- CP-element group 4: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_Update/cca
      -- 
    cca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_258_call_ack_1, ack => getQueuePointer_CP_134_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_sample_start_
      -- CP-element group 5: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Sample/crr
      -- 
    crr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(5), ack => call_stmt_267_call_req_0); -- 
    getQueuePointer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "getQueuePointer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getQueuePointer_CP_134_elements(2) & getQueuePointer_CP_134_elements(11);
      gj_getQueuePointer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getQueuePointer_CP_134_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_sample_completed_
      -- CP-element group 6: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Sample/cra
      -- 
    cra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_267_call_ack_0, ack => getQueuePointer_CP_134_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_update_completed_
      -- CP-element group 7: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Update/$exit
      -- CP-element group 7: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_267_Update/cca
      -- 
    cca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_267_call_ack_1, ack => getQueuePointer_CP_134_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_sample_start_
      -- CP-element group 8: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Sample/rr
      -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointer_CP_134_elements(8), ack => CONCAT_u32_u64_271_inst_req_0); -- 
    getQueuePointer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "getQueuePointer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getQueuePointer_CP_134_elements(4) & getQueuePointer_CP_134_elements(7);
      gj_getQueuePointer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getQueuePointer_CP_134_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_sample_completed_
      -- CP-element group 9: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Sample/ra
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_271_inst_ack_0, ack => getQueuePointer_CP_134_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 $exit
      -- CP-element group 10: 	 assign_stmt_251_to_assign_stmt_272/$exit
      -- CP-element group 10: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_update_completed_
      -- CP-element group 10: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Update/$exit
      -- CP-element group 10: 	 assign_stmt_251_to_assign_stmt_272/CONCAT_u32_u64_271_Update/ca
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_271_inst_ack_1, ack => getQueuePointer_CP_134_elements(10)); -- 
    -- CP-element group 11:  transition  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	4 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 assign_stmt_251_to_assign_stmt_272/call_stmt_258_call_stmt_267_delay
      -- 
    -- Element group getQueuePointer_CP_134_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => getQueuePointer_CP_134_elements(4), ack => getQueuePointer_CP_134_elements(11), clk => clk, reset =>reset);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_263_wire : std_logic_vector(7 downto 0);
    signal R_READMEM_252_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_259_wire_constant : std_logic_vector(0 downto 0);
    signal base_idx_251 : std_logic_vector(7 downto 0);
    signal call_getBaseIndex_expr_250_wire : std_logic_vector(7 downto 0);
    signal konst_253_wire_constant : std_logic_vector(3 downto 0);
    signal konst_260_wire_constant : std_logic_vector(3 downto 0);
    signal konst_262_wire_constant : std_logic_vector(7 downto 0);
    signal qptr_h_258 : std_logic_vector(31 downto 0);
    signal qptr_l_267 : std_logic_vector(31 downto 0);
    signal type_cast_256_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_265_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_252_wire_constant <= "1";
    R_READMEM_259_wire_constant <= "1";
    konst_253_wire_constant <= "1111";
    konst_260_wire_constant <= "1111";
    konst_262_wire_constant <= "00000001";
    type_cast_256_wire_constant <= "00000000000000000000000000000000";
    type_cast_265_wire_constant <= "00000000000000000000000000000000";
    W_base_idx_247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_base_idx_247_inst_req_0;
      W_base_idx_247_inst_ack_0<= wack(0);
      rreq(0) <= W_base_idx_247_inst_req_1;
      W_base_idx_247_inst_ack_1<= rack(0);
      W_base_idx_247_inst : InterlockBuffer generic map ( -- 
        name => "W_base_idx_247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_getBaseIndex_expr_250_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => base_idx_251,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- flow through binary operator ADD_u8_u8_263_inst
    ADD_u8_u8_263_wire <= std_logic_vector(unsigned(base_idx_251) + unsigned(konst_262_wire_constant));
    -- shared split operator group (1) : CONCAT_u32_u64_271_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= qptr_h_258 & qptr_l_267;
      qptr_buffer <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_271_inst_req_0;
      CONCAT_u32_u64_271_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_271_inst_req_1;
      CONCAT_u32_u64_271_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    volatile_operator_getBaseIndex_450: getBaseIndex_Volatile port map(queue_type => queue_type_buffer, server_id => server_id_buffer, base_index => call_getBaseIndex_expr_250_wire); 
    -- shared call operator group (1) : call_stmt_258_call call_stmt_267_call 
    accessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_258_call_req_0;
      reqL_unguarded(0) <= call_stmt_267_call_req_0;
      call_stmt_258_call_ack_0 <= ackL_unguarded(1);
      call_stmt_267_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_258_call_req_1;
      reqR_unguarded(0) <= call_stmt_267_call_req_1;
      call_stmt_258_call_ack_1 <= ackR_unguarded(1);
      call_stmt_267_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessRegister_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "accessRegister_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "accessRegister_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_READMEM_252_wire_constant & konst_253_wire_constant & base_idx_251 & type_cast_256_wire_constant & R_READMEM_259_wire_constant & konst_260_wire_constant & ADD_u8_u8_263_wire & type_cast_265_wire_constant;
      qptr_h_258 <= data_out(63 downto 32);
      qptr_l_267 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 90,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getQueuePointer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    q_base_address : in  std_logic_vector(63 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
    accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
    accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
    accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
    accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
    accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(63 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_1302_start: Boolean;
  signal getQueuePointers_CP_1302_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueReadIndex is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessQueueWriteIndex is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_979_call_req_0 : boolean;
  signal call_stmt_979_call_ack_0 : boolean;
  signal call_stmt_979_call_req_1 : boolean;
  signal call_stmt_979_call_ack_1 : boolean;
  signal call_stmt_986_call_req_0 : boolean;
  signal call_stmt_986_call_ack_0 : boolean;
  signal call_stmt_986_call_req_1 : boolean;
  signal call_stmt_986_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_1302_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_1302_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_1302_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_1302_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_1302: Block -- control-path 
    signal getQueuePointers_CP_1302_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_1302_elements(0) <= getQueuePointers_CP_1302_start;
    getQueuePointers_CP_1302_symbol <= getQueuePointers_CP_1302_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/$entry
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_sample_start_
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_update_start_
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Sample/$entry
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Sample/crr
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Update/$entry
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Update/ccr
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_update_start_
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Update/$entry
      -- CP-element group 0: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Update/ccr
      -- 
    ccr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1302_elements(0), ack => call_stmt_986_call_req_1); -- 
    crr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1302_elements(0), ack => call_stmt_979_call_req_0); -- 
    ccr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1302_elements(0), ack => call_stmt_979_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_sample_completed_
      -- CP-element group 1: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Sample/$exit
      -- CP-element group 1: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Sample/cra
      -- 
    cra_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_979_call_ack_0, ack => getQueuePointers_CP_1302_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_update_completed_
      -- CP-element group 2: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Update/$exit
      -- CP-element group 2: 	 call_stmt_979_to_call_stmt_986/call_stmt_979_Update/cca
      -- CP-element group 2: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_sample_start_
      -- CP-element group 2: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Sample/$entry
      -- CP-element group 2: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Sample/crr
      -- 
    cca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_979_call_ack_1, ack => getQueuePointers_CP_1302_elements(2)); -- 
    crr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1302_elements(2), ack => call_stmt_986_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_sample_completed_
      -- CP-element group 3: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Sample/$exit
      -- CP-element group 3: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Sample/cra
      -- 
    cra_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_986_call_ack_0, ack => getQueuePointers_CP_1302_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_979_to_call_stmt_986/$exit
      -- CP-element group 4: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_update_completed_
      -- CP-element group 4: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Update/$exit
      -- CP-element group 4: 	 call_stmt_979_to_call_stmt_986/call_stmt_986_Update/cca
      -- 
    cca_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_986_call_ack_1, ack => getQueuePointers_CP_1302_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_READMEM_974_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_981_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_984_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_974_wire_constant <= "1";
    R_READMEM_981_wire_constant <= "1";
    type_cast_977_wire_constant <= "00000000000000000000000000000000";
    type_cast_984_wire_constant <= "00000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_979_call 
    accessQueueReadIndex_call_group_0: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_979_call_req_0;
      call_stmt_979_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_979_call_req_1;
      call_stmt_979_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueReadIndex_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueReadIndex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_974_wire_constant & q_base_address_buffer & type_cast_977_wire_constant;
      rp_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueReadIndex_call_reqs(0),
          ackR => accessQueueReadIndex_call_acks(0),
          dataR => accessQueueReadIndex_call_data(104 downto 0),
          tagR => accessQueueReadIndex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueReadIndex_return_acks(0), -- cross-over
          ackL => accessQueueReadIndex_return_reqs(0), -- cross-over
          dataL => accessQueueReadIndex_return_data(31 downto 0),
          tagL => accessQueueReadIndex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_986_call 
    accessQueueWriteIndex_call_group_1: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_986_call_req_0;
      call_stmt_986_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_986_call_req_1;
      call_stmt_986_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueWriteIndex_call_group_1_gI: SplitGuardInterface generic map(name => "accessQueueWriteIndex_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_981_wire_constant & q_base_address_buffer & type_cast_984_wire_constant;
      wp_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueWriteIndex_call_reqs(0),
          ackR => accessQueueWriteIndex_call_acks(0),
          dataR => accessQueueWriteIndex_call_data(104 downto 0),
          tagR => accessQueueWriteIndex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueWriteIndex_return_acks(0), -- cross-over
          ackL => accessQueueWriteIndex_return_reqs(0), -- cross-over
          dataL => accessQueueWriteIndex_return_data(31 downto 0),
          tagL => accessQueueWriteIndex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    q_base_address : in  std_logic_vector(63 downto 0);
    total_msgs : out  std_logic_vector(31 downto 0);
    accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
    accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
    accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTotalMessages;
architecture getTotalMessages_arch of getTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(63 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal total_msgs_update_enable: Boolean;
  signal getTotalMessages_CP_1396_start: Boolean;
  signal getTotalMessages_CP_1396_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueTotalMsgs is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1038_call_req_0 : boolean;
  signal call_stmt_1038_call_ack_0 : boolean;
  signal call_stmt_1038_call_req_1 : boolean;
  signal call_stmt_1038_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTotalMessages_CP_1396_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= total_msgs_buffer;
  total_msgs <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_1396_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTotalMessages_CP_1396_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_1396_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTotalMessages_CP_1396: Block -- control-path 
    signal getTotalMessages_CP_1396_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    getTotalMessages_CP_1396_elements(0) <= getTotalMessages_CP_1396_start;
    getTotalMessages_CP_1396_symbol <= getTotalMessages_CP_1396_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1038/$entry
      -- CP-element group 0: 	 call_stmt_1038/call_stmt_1038_sample_start_
      -- CP-element group 0: 	 call_stmt_1038/call_stmt_1038_update_start_
      -- CP-element group 0: 	 call_stmt_1038/call_stmt_1038_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1038/call_stmt_1038_Sample/crr
      -- CP-element group 0: 	 call_stmt_1038/call_stmt_1038_Update/$entry
      -- CP-element group 0: 	 call_stmt_1038/call_stmt_1038_Update/ccr
      -- 
    crr_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_1396_elements(0), ack => call_stmt_1038_call_req_0); -- 
    ccr_1414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_1396_elements(0), ack => call_stmt_1038_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1038/call_stmt_1038_sample_completed_
      -- CP-element group 1: 	 call_stmt_1038/call_stmt_1038_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1038/call_stmt_1038_Sample/cra
      -- 
    cra_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1038_call_ack_0, ack => getTotalMessages_CP_1396_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1038/$exit
      -- CP-element group 2: 	 call_stmt_1038/call_stmt_1038_update_completed_
      -- CP-element group 2: 	 call_stmt_1038/call_stmt_1038_Update/$exit
      -- CP-element group 2: 	 call_stmt_1038/call_stmt_1038_Update/cca
      -- 
    cca_1415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1038_call_ack_1, ack => getTotalMessages_CP_1396_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_READMEM_1033_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_1033_wire_constant <= "1";
    type_cast_1036_wire_constant <= "00000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_1038_call 
    accessQueueTotalMsgs_call_group_0: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1038_call_req_0;
      call_stmt_1038_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1038_call_req_1;
      call_stmt_1038_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueTotalMsgs_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueTotalMsgs_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_1033_wire_constant & q_base_address_buffer & type_cast_1036_wire_constant;
      total_msgs_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueTotalMsgs_call_reqs(0),
          ackR => accessQueueTotalMsgs_call_acks(0),
          dataR => accessQueueTotalMsgs_call_data(104 downto 0),
          tagR => accessQueueTotalMsgs_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueTotalMsgs_return_acks(0), -- cross-over
          ackL => accessQueueTotalMsgs_return_reqs(0), -- cross-over
          dataL => accessQueueTotalMsgs_return_data(31 downto 0),
          tagL => accessQueueTotalMsgs_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    server_index : in  std_logic_vector(7 downto 0);
    pkt_pointer : out  std_logic_vector(63 downto 0);
    status : out  std_logic_vector(0 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(17 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(64 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 65)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal server_index_buffer :  std_logic_vector(7 downto 0);
  signal server_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(63 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_3989_start: Boolean;
  signal getTxPacketPointerFromServer_CP_3989_symbol: Boolean;
  -- volatile/operator module components. 
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_r_data : out  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueMisc_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueMisc_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueMisc_call_data : out  std_logic_vector(104 downto 0);
      accessQueueMisc_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueMisc_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueMisc_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueMisc_return_data : in   std_logic_vector(31 downto 0);
      accessQueueMisc_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(103 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(63 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_2136_call_req_0 : boolean;
  signal call_stmt_2136_call_ack_0 : boolean;
  signal call_stmt_2136_call_req_1 : boolean;
  signal call_stmt_2136_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 16) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(15 downto 8) <= server_index;
  server_index_buffer <= in_buffer_data_out(15 downto 8);
  in_buffer_data_in(tag_length + 15 downto 16) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 15 downto 16);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 1,3 => 7);
    constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 7);
    constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 4); -- 
  begin -- 
    preds <= tag_update_enable & server_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_3989_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 65) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(64 downto 64) <= status_buffer;
  status <= out_buffer_data_out(64 downto 64);
  out_buffer_data_in(tag_length + 64 downto 65) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 64 downto 65);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_3989_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_3989_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_3989_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_3989: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_3989_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_3989_elements(0) <= getTxPacketPointerFromServer_CP_3989_start;
    getTxPacketPointerFromServer_CP_3989_symbol <= getTxPacketPointerFromServer_CP_3989_elements(14);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_2136/$entry
      -- 
    getTxPacketPointerFromServer_CP_3989_elements(1) <= getTxPacketPointerFromServer_CP_3989_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	10 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_2136/tag_update_enable
      -- CP-element group 2: 	 call_stmt_2136/tag_update_enable_out
      -- 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_3989_elements(8);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3989_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	8 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	11 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_2136/server_index_update_enable
      -- CP-element group 3: 	 call_stmt_2136/server_index_update_enable_out
      -- 
    getTxPacketPointerFromServer_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_3989_elements(8);
      gj_getTxPacketPointerFromServer_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3989_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	12 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_2136/pkt_pointer_update_enable
      -- CP-element group 4: 	 call_stmt_2136/pkt_pointer_update_enable_in
      -- 
    getTxPacketPointerFromServer_CP_3989_elements(4) <= getTxPacketPointerFromServer_CP_3989_elements(12);
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	13 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_2136/status_update_enable
      -- CP-element group 5: 	 call_stmt_2136/status_update_enable_in
      -- 
    getTxPacketPointerFromServer_CP_3989_elements(5) <= getTxPacketPointerFromServer_CP_3989_elements(13);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_2136/call_stmt_2136_sample_start_
      -- CP-element group 6: 	 call_stmt_2136/call_stmt_2136_Sample/$entry
      -- CP-element group 6: 	 call_stmt_2136/call_stmt_2136_Sample/crr
      -- 
    crr_4010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_3989_elements(6), ack => call_stmt_2136_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_3989_elements(1) & getTxPacketPointerFromServer_CP_3989_elements(8);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3989_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	5 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_2136/call_stmt_2136_update_start_
      -- CP-element group 7: 	 call_stmt_2136/call_stmt_2136_Update/$entry
      -- CP-element group 7: 	 call_stmt_2136/call_stmt_2136_Update/ccr
      -- 
    ccr_4015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_3989_elements(7), ack => call_stmt_2136_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_3989_elements(4) & getTxPacketPointerFromServer_CP_3989_elements(5) & getTxPacketPointerFromServer_CP_3989_elements(9);
      gj_getTxPacketPointerFromServer_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3989_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_2136/call_stmt_2136_sample_completed_
      -- CP-element group 8: 	 call_stmt_2136/call_stmt_2136_Sample/$exit
      -- CP-element group 8: 	 call_stmt_2136/call_stmt_2136_Sample/cra
      -- 
    cra_4011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2136_call_ack_0, ack => getTxPacketPointerFromServer_CP_3989_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 call_stmt_2136/$exit
      -- CP-element group 9: 	 call_stmt_2136/call_stmt_2136_update_completed_
      -- CP-element group 9: 	 call_stmt_2136/call_stmt_2136_Update/$exit
      -- CP-element group 9: 	 call_stmt_2136/call_stmt_2136_Update/cca
      -- 
    cca_4016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2136_call_ack_1, ack => getTxPacketPointerFromServer_CP_3989_elements(9)); -- 
    -- CP-element group 10:  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 tag_update_enable
      -- 
    getTxPacketPointerFromServer_CP_3989_elements(10) <= getTxPacketPointerFromServer_CP_3989_elements(2);
    -- CP-element group 11:  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	3 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 server_index_update_enable
      -- 
    getTxPacketPointerFromServer_CP_3989_elements(11) <= getTxPacketPointerFromServer_CP_3989_elements(3);
    -- CP-element group 12:  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	4 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 pkt_pointer_update_enable
      -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	5 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 status_update_enable
      -- 
    -- CP-element group 14:  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 $exit
      -- 
    getTxPacketPointerFromServer_CP_3989_elements(14) <= getTxPacketPointerFromServer_CP_3989_elements(9);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_3989_elements(12) <= pkt_pointer_update_enable;
    getTxPacketPointerFromServer_CP_3989_elements(13) <= status_update_enable;
    -- hookup: output from control-path 
    tag_update_enable <= getTxPacketPointerFromServer_CP_3989_elements(10);
    server_index_update_enable <= getTxPacketPointerFromServer_CP_3989_elements(11);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_TXQUEUE_2132_wire_constant : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    R_TXQUEUE_2132_wire_constant <= "01";
    -- shared call operator group (0) : call_stmt_2136_call 
    popFromQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2136_call_req_0;
      call_stmt_2136_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2136_call_req_1;
      call_stmt_2136_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_0_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_TXQUEUE_2132_wire_constant & server_index_buffer;
      pkt_pointer_buffer <= data_out(64 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 18,
        owidth => 18,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(17 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 65,
          owidth => 65,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(64 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity incrementNumberOfPacketsReceived is -- 
  generic (tag_length : integer); 
  port ( -- 
    incrementRegister_call_reqs : out  std_logic_vector(0 downto 0);
    incrementRegister_call_acks : in   std_logic_vector(0 downto 0);
    incrementRegister_call_data : out  std_logic_vector(7 downto 0);
    incrementRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    incrementRegister_return_reqs : out  std_logic_vector(0 downto 0);
    incrementRegister_return_acks : in   std_logic_vector(0 downto 0);
    incrementRegister_return_data : in   std_logic_vector(31 downto 0);
    incrementRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity incrementNumberOfPacketsReceived;
architecture incrementNumberOfPacketsReceived_arch of incrementNumberOfPacketsReceived is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal incrementNumberOfPacketsReceived_CP_2687_start: Boolean;
  signal incrementNumberOfPacketsReceived_CP_2687_symbol: Boolean;
  -- volatile/operator module components. 
  component incrementRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      reg_index : in  std_logic_vector(7 downto 0);
      incremented_value : out  std_logic_vector(31 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1720_call_ack_1 : boolean;
  signal call_stmt_1720_call_req_1 : boolean;
  signal call_stmt_1720_call_ack_0 : boolean;
  signal call_stmt_1720_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "incrementNumberOfPacketsReceived_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  incrementNumberOfPacketsReceived_CP_2687_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "incrementNumberOfPacketsReceived_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= incrementNumberOfPacketsReceived_CP_2687_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= incrementNumberOfPacketsReceived_CP_2687_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= incrementNumberOfPacketsReceived_CP_2687_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  incrementNumberOfPacketsReceived_CP_2687: Block -- control-path 
    signal incrementNumberOfPacketsReceived_CP_2687_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    incrementNumberOfPacketsReceived_CP_2687_elements(0) <= incrementNumberOfPacketsReceived_CP_2687_start;
    incrementNumberOfPacketsReceived_CP_2687_symbol <= incrementNumberOfPacketsReceived_CP_2687_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_1720/call_stmt_1720_update_start_
      -- CP-element group 0: 	 call_stmt_1720/call_stmt_1720_sample_start_
      -- CP-element group 0: 	 call_stmt_1720/$entry
      -- CP-element group 0: 	 call_stmt_1720/call_stmt_1720_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1720/call_stmt_1720_Update/ccr
      -- CP-element group 0: 	 call_stmt_1720/call_stmt_1720_Update/$entry
      -- CP-element group 0: 	 call_stmt_1720/call_stmt_1720_Sample/crr
      -- 
    crr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementNumberOfPacketsReceived_CP_2687_elements(0), ack => call_stmt_1720_call_req_0); -- 
    ccr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementNumberOfPacketsReceived_CP_2687_elements(0), ack => call_stmt_1720_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1720/call_stmt_1720_sample_completed_
      -- CP-element group 1: 	 call_stmt_1720/call_stmt_1720_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1720/call_stmt_1720_Sample/cra
      -- 
    cra_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1720_call_ack_0, ack => incrementNumberOfPacketsReceived_CP_2687_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_1720/$exit
      -- CP-element group 2: 	 call_stmt_1720/call_stmt_1720_update_completed_
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1720/call_stmt_1720_Update/cca
      -- CP-element group 2: 	 call_stmt_1720/call_stmt_1720_Update/$exit
      -- 
    cca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1720_call_ack_1, ack => incrementNumberOfPacketsReceived_CP_2687_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ignore_val_1720 : std_logic_vector(31 downto 0);
    signal konst_1718_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1718_wire_constant <= "11010011";
    -- shared call operator group (0) : call_stmt_1720_call 
    incrementRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1720_call_req_0;
      call_stmt_1720_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1720_call_req_1;
      call_stmt_1720_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      incrementRegister_call_group_0_gI: SplitGuardInterface generic map(name => "incrementRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_1718_wire_constant;
      ignore_val_1720 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 8,
        owidth => 8,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => incrementRegister_call_reqs(0),
          ackR => incrementRegister_call_acks(0),
          dataR => incrementRegister_call_data(7 downto 0),
          tagR => incrementRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => incrementRegister_return_acks(0), -- cross-over
          ackL => incrementRegister_return_reqs(0), -- cross-over
          dataL => incrementRegister_return_data(31 downto 0),
          tagL => incrementRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end incrementNumberOfPacketsReceived_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity incrementNumberOfPacketsTransmitted is -- 
  generic (tag_length : integer); 
  port ( -- 
    incrementRegister_call_reqs : out  std_logic_vector(0 downto 0);
    incrementRegister_call_acks : in   std_logic_vector(0 downto 0);
    incrementRegister_call_data : out  std_logic_vector(7 downto 0);
    incrementRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    incrementRegister_return_reqs : out  std_logic_vector(0 downto 0);
    incrementRegister_return_acks : in   std_logic_vector(0 downto 0);
    incrementRegister_return_data : in   std_logic_vector(31 downto 0);
    incrementRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity incrementNumberOfPacketsTransmitted;
architecture incrementNumberOfPacketsTransmitted_arch of incrementNumberOfPacketsTransmitted is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal incrementNumberOfPacketsTransmitted_CP_4024_start: Boolean;
  signal incrementNumberOfPacketsTransmitted_CP_4024_symbol: Boolean;
  -- volatile/operator module components. 
  component incrementRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      reg_index : in  std_logic_vector(7 downto 0);
      incremented_value : out  std_logic_vector(31 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_2144_call_req_0 : boolean;
  signal call_stmt_2144_call_ack_0 : boolean;
  signal call_stmt_2144_call_req_1 : boolean;
  signal call_stmt_2144_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "incrementNumberOfPacketsTransmitted_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  incrementNumberOfPacketsTransmitted_CP_4024_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "incrementNumberOfPacketsTransmitted_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= incrementNumberOfPacketsTransmitted_CP_4024_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= incrementNumberOfPacketsTransmitted_CP_4024_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= incrementNumberOfPacketsTransmitted_CP_4024_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  incrementNumberOfPacketsTransmitted_CP_4024: Block -- control-path 
    signal incrementNumberOfPacketsTransmitted_CP_4024_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    incrementNumberOfPacketsTransmitted_CP_4024_elements(0) <= incrementNumberOfPacketsTransmitted_CP_4024_start;
    incrementNumberOfPacketsTransmitted_CP_4024_symbol <= incrementNumberOfPacketsTransmitted_CP_4024_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_2144/$entry
      -- CP-element group 0: 	 call_stmt_2144/call_stmt_2144_sample_start_
      -- CP-element group 0: 	 call_stmt_2144/call_stmt_2144_update_start_
      -- CP-element group 0: 	 call_stmt_2144/call_stmt_2144_Sample/$entry
      -- CP-element group 0: 	 call_stmt_2144/call_stmt_2144_Sample/crr
      -- CP-element group 0: 	 call_stmt_2144/call_stmt_2144_Update/$entry
      -- CP-element group 0: 	 call_stmt_2144/call_stmt_2144_Update/ccr
      -- 
    crr_4037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementNumberOfPacketsTransmitted_CP_4024_elements(0), ack => call_stmt_2144_call_req_0); -- 
    ccr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementNumberOfPacketsTransmitted_CP_4024_elements(0), ack => call_stmt_2144_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_2144/call_stmt_2144_sample_completed_
      -- CP-element group 1: 	 call_stmt_2144/call_stmt_2144_Sample/$exit
      -- CP-element group 1: 	 call_stmt_2144/call_stmt_2144_Sample/cra
      -- 
    cra_4038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2144_call_ack_0, ack => incrementNumberOfPacketsTransmitted_CP_4024_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_2144/$exit
      -- CP-element group 2: 	 call_stmt_2144/call_stmt_2144_update_completed_
      -- CP-element group 2: 	 call_stmt_2144/call_stmt_2144_Update/$exit
      -- CP-element group 2: 	 call_stmt_2144/call_stmt_2144_Update/cca
      -- 
    cca_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2144_call_ack_1, ack => incrementNumberOfPacketsTransmitted_CP_4024_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ignore_val_2144 : std_logic_vector(31 downto 0);
    signal konst_2142_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_2142_wire_constant <= "11010010";
    -- shared call operator group (0) : call_stmt_2144_call 
    incrementRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2144_call_req_0;
      call_stmt_2144_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2144_call_req_1;
      call_stmt_2144_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      incrementRegister_call_group_0_gI: SplitGuardInterface generic map(name => "incrementRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_2142_wire_constant;
      ignore_val_2144 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 8,
        owidth => 8,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => incrementRegister_call_reqs(0),
          ackR => incrementRegister_call_acks(0),
          dataR => incrementRegister_call_data(7 downto 0),
          tagR => incrementRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => incrementRegister_return_acks(0), -- cross-over
          ackL => incrementRegister_return_reqs(0), -- cross-over
          dataL => incrementRegister_return_data(31 downto 0),
          tagL => incrementRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end incrementNumberOfPacketsTransmitted_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity incrementRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    reg_index : in  std_logic_vector(7 downto 0);
    incremented_value : out  std_logic_vector(31 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_call_acks : in   std_logic_vector(0 downto 0);
    accessRegister_call_data : out  std_logic_vector(44 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_return_acks : in   std_logic_vector(0 downto 0);
    accessRegister_return_data : in   std_logic_vector(31 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity incrementRegister;
architecture incrementRegister_arch of incrementRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal reg_index_buffer :  std_logic_vector(7 downto 0);
  signal reg_index_update_enable: Boolean;
  -- output port buffer signals
  signal incremented_value_buffer :  std_logic_vector(31 downto 0);
  signal incremented_value_update_enable: Boolean;
  signal incrementRegister_CP_2652_start: Boolean;
  signal incrementRegister_CP_2652_symbol: Boolean;
  -- volatile/operator module components. 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1703_call_req_0 : boolean;
  signal call_stmt_1715_call_ack_1 : boolean;
  signal call_stmt_1715_call_req_1 : boolean;
  signal call_stmt_1715_call_ack_0 : boolean;
  signal call_stmt_1715_call_req_0 : boolean;
  signal call_stmt_1703_call_ack_1 : boolean;
  signal call_stmt_1703_call_req_1 : boolean;
  signal call_stmt_1703_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "incrementRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 8) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= reg_index;
  reg_index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(tag_length + 7 downto 8) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 7 downto 8);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  incrementRegister_CP_2652_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "incrementRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= incremented_value_buffer;
  incremented_value <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= incrementRegister_CP_2652_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= incrementRegister_CP_2652_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= incrementRegister_CP_2652_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  incrementRegister_CP_2652: Block -- control-path 
    signal incrementRegister_CP_2652_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    incrementRegister_CP_2652_elements(0) <= incrementRegister_CP_2652_start;
    incrementRegister_CP_2652_symbol <= incrementRegister_CP_2652_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_sample_start_
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Sample/crr
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/$entry
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Update/ccr
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Update/$entry
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Update/ccr
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Update/$entry
      -- CP-element group 0: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_update_start_
      -- 
    crr_2665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementRegister_CP_2652_elements(0), ack => call_stmt_1703_call_req_0); -- 
    ccr_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementRegister_CP_2652_elements(0), ack => call_stmt_1703_call_req_1); -- 
    ccr_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementRegister_CP_2652_elements(0), ack => call_stmt_1715_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Sample/cra
      -- CP-element group 1: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_sample_completed_
      -- 
    cra_2666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1703_call_ack_0, ack => incrementRegister_CP_2652_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_update_completed_
      -- CP-element group 2: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Update/cca
      -- CP-element group 2: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_Update/$exit
      -- 
    cca_2671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1703_call_ack_1, ack => incrementRegister_CP_2652_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	5 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Sample/cra
      -- CP-element group 3: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_sample_completed_
      -- 
    cra_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1715_call_ack_0, ack => incrementRegister_CP_2652_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 call_stmt_1703_to_call_stmt_1715/$exit
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Update/cca
      -- CP-element group 4: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Update/$exit
      -- CP-element group 4: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_update_completed_
      -- 
    cca_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1715_call_ack_1, ack => incrementRegister_CP_2652_elements(4)); -- 
    -- CP-element group 5:  transition  output  delay-element  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	3 
    -- CP-element group 5:  members (4) 
      -- CP-element group 5: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1703_call_stmt_1715_delay
      -- CP-element group 5: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Sample/crr
      -- CP-element group 5: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_Sample/$entry
      -- CP-element group 5: 	 call_stmt_1703_to_call_stmt_1715/call_stmt_1715_sample_start_
      -- 
    crr_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => incrementRegister_CP_2652_elements(5), ack => call_stmt_1715_call_req_0); -- 
    -- Element group incrementRegister_CP_2652_elements(5) is a control-delay.
    cp_element_5_delay: control_delay_element  generic map(name => " 5_delay", delay_value => 1)  port map(req => incrementRegister_CP_2652_elements(2), ack => incrementRegister_CP_2652_elements(5), clk => clk, reset =>reset);
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_1698_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1706_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1711_wire_constant : std_logic_vector(3 downto 0);
    signal rval_1703 : std_logic_vector(31 downto 0);
    signal rval_ignore_1715 : std_logic_vector(31 downto 0);
    signal type_cast_1697_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1710_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1698_wire_constant <= "1111";
    konst_1706_wire_constant <= "00000000000000000000000000000001";
    konst_1711_wire_constant <= "1111";
    type_cast_1697_wire_constant <= "1";
    type_cast_1701_wire_constant <= "00000000000000000000000000000000";
    type_cast_1710_wire_constant <= "0";
    -- flow through binary operator ADD_u32_u32_1707_inst
    incremented_value_buffer <= std_logic_vector(unsigned(rval_1703) + unsigned(konst_1706_wire_constant));
    -- shared call operator group (0) : call_stmt_1703_call call_stmt_1715_call 
    accessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1703_call_req_0;
      reqL_unguarded(0) <= call_stmt_1715_call_req_0;
      call_stmt_1703_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1715_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1703_call_req_1;
      reqR_unguarded(0) <= call_stmt_1715_call_req_1;
      call_stmt_1703_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1715_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1697_wire_constant & konst_1698_wire_constant & reg_index_buffer & type_cast_1701_wire_constant & type_cast_1710_wire_constant & konst_1711_wire_constant & reg_index_buffer & incremented_value_buffer;
      rval_1703 <= data_out(63 downto 32);
      rval_ignore_1715 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 90,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end incrementRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    max_addr_offset : in  std_logic_vector(15 downto 0);
    rx_buffer_pointer : in  std_logic_vector(63 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(71 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(15 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(103 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(106 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 88)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal max_addr_offset_buffer :  std_logic_vector(15 downto 0);
  signal max_addr_offset_update_enable: Boolean;
  signal rx_buffer_pointer_buffer :  std_logic_vector(63 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_2250_start: Boolean;
  signal loadBuffer_CP_2250_symbol: Boolean;
  -- volatile/operator module components. 
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      buf_pointer : in  std_logic_vector(63 downto 0);
      addr_offset : out  std_logic_vector(15 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      max_addr_offset : in  std_logic_vector(15 downto 0);
      base_buf_pointer : in  std_logic_vector(63 downto 0);
      addr_offset : in  std_logic_vector(15 downto 0);
      packet_size_11 : out  std_logic_vector(10 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      base_buffer_pointer : in  std_logic_vector(63 downto 0);
      max_addr_offset : in  std_logic_vector(15 downto 0);
      packet_size : in  std_logic_vector(10 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1559_call_ack_1 : boolean;
  signal W_bad_packet_identifier_1462_delayed_8_0_1541_inst_ack_1 : boolean;
  signal call_stmt_1559_call_req_1 : boolean;
  signal W_tag_1463_delayed_8_0_1544_inst_req_0 : boolean;
  signal W_tag_1463_delayed_8_0_1544_inst_ack_0 : boolean;
  signal W_tag_1463_delayed_8_0_1544_inst_req_1 : boolean;
  signal W_max_addr_offset_1455_delayed_4_0_1527_inst_req_0 : boolean;
  signal W_max_addr_offset_1455_delayed_4_0_1527_inst_ack_0 : boolean;
  signal W_tag_1463_delayed_8_0_1544_inst_ack_1 : boolean;
  signal call_stmt_1522_call_req_0 : boolean;
  signal W_max_addr_offset_1455_delayed_4_0_1527_inst_req_1 : boolean;
  signal W_max_addr_offset_1455_delayed_4_0_1527_inst_ack_1 : boolean;
  signal call_stmt_1522_call_ack_0 : boolean;
  signal W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_ack_1 : boolean;
  signal call_stmt_1522_call_req_1 : boolean;
  signal call_stmt_1522_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_ack_0 : boolean;
  signal W_bad_packet_identifier_1462_delayed_8_0_1541_inst_req_1 : boolean;
  signal W_bad_packet_identifier_1462_delayed_8_0_1541_inst_ack_0 : boolean;
  signal W_bad_packet_identifier_1462_delayed_8_0_1541_inst_req_0 : boolean;
  signal call_stmt_1559_call_ack_0 : boolean;
  signal call_stmt_1559_call_req_0 : boolean;
  signal W_max_addr_offset_1465_delayed_8_0_1550_inst_ack_1 : boolean;
  signal W_max_addr_offset_1465_delayed_8_0_1550_inst_req_1 : boolean;
  signal W_tag_1454_delayed_4_0_1524_inst_ack_1 : boolean;
  signal W_tag_1454_delayed_4_0_1524_inst_req_1 : boolean;
  signal W_tag_1454_delayed_4_0_1524_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_ack_1 : boolean;
  signal W_tag_1454_delayed_4_0_1524_inst_req_0 : boolean;
  signal W_max_addr_offset_1465_delayed_8_0_1550_inst_ack_0 : boolean;
  signal call_stmt_1540_call_ack_1 : boolean;
  signal call_stmt_1540_call_req_1 : boolean;
  signal call_stmt_1540_call_ack_0 : boolean;
  signal W_max_addr_offset_1465_delayed_8_0_1550_inst_req_0 : boolean;
  signal call_stmt_1540_call_req_0 : boolean;
  signal W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 88) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(23 downto 8) <= max_addr_offset;
  max_addr_offset_buffer <= in_buffer_data_out(23 downto 8);
  in_buffer_data_in(87 downto 24) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(87 downto 24);
  in_buffer_data_in(tag_length + 87 downto 88) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 87 downto 88);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 31);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 31);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= tag_update_enable & max_addr_offset_update_enable & rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_2250_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_2250_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_2250_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_2250_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_2250: Block -- control-path 
    signal loadBuffer_CP_2250_elements: BooleanArray(50 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_2250_elements(0) <= loadBuffer_CP_2250_start;
    loadBuffer_CP_2250_symbol <= loadBuffer_CP_2250_elements(50);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	34 
    -- CP-element group 1: 	38 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1522_to_call_stmt_1559/$entry
      -- 
    loadBuffer_CP_2250_elements(1) <= loadBuffer_CP_2250_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	32 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	46 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1522_to_call_stmt_1559/tag_update_enable_out
      -- CP-element group 2: 	 call_stmt_1522_to_call_stmt_1559/tag_update_enable
      -- 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(8) & loadBuffer_CP_2250_elements(12) & loadBuffer_CP_2250_elements(32);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	16 
    -- CP-element group 3: 	40 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	47 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1522_to_call_stmt_1559/max_addr_offset_update_enable_out
      -- CP-element group 3: 	 call_stmt_1522_to_call_stmt_1559/max_addr_offset_update_enable
      -- 
    loadBuffer_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(16) & loadBuffer_CP_2250_elements(40);
      gj_loadBuffer_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	20 
    -- CP-element group 4: 	36 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	48 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 call_stmt_1522_to_call_stmt_1559/rx_buffer_pointer_update_enable_out
      -- CP-element group 4: 	 call_stmt_1522_to_call_stmt_1559/rx_buffer_pointer_update_enable
      -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(8) & loadBuffer_CP_2250_elements(20) & loadBuffer_CP_2250_elements(36);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	49 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	23 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 call_stmt_1522_to_call_stmt_1559/bad_packet_identifier_update_enable_in
      -- CP-element group 5: 	 call_stmt_1522_to_call_stmt_1559/bad_packet_identifier_update_enable
      -- 
    loadBuffer_CP_2250_elements(5) <= loadBuffer_CP_2250_elements(49);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	45 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_sample_start_
      -- CP-element group 6: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Sample/crr
      -- 
    crr_2271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(6), ack => call_stmt_1522_call_req_0); -- 
    loadBuffer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(8) & loadBuffer_CP_2250_elements(45);
      gj_loadBuffer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: 	24 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_update_start_
      -- CP-element group 7: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Update/$entry
      -- CP-element group 7: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Update/ccr
      -- 
    ccr_2276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(7), ack => call_stmt_1522_call_req_1); -- 
    loadBuffer_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(24);
      gj_loadBuffer_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_sample_completed_
      -- CP-element group 8: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Sample/$exit
      -- CP-element group 8: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Sample/cra
      -- 
    cra_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1522_call_ack_0, ack => loadBuffer_CP_2250_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	18 
    -- CP-element group 9: 	22 
    -- CP-element group 9: 	26 
    -- CP-element group 9: 	30 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	38 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_update_completed_
      -- CP-element group 9: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Update/$exit
      -- CP-element group 9: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1522_Update/cca
      -- CP-element group 9: 	 call_stmt_1522_to_call_stmt_1559/barrier_stmt_1523_update_completed_
      -- 
    cca_2277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1522_call_ack_1, ack => loadBuffer_CP_2250_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_sample_start_
      -- CP-element group 10: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Sample/req
      -- CP-element group 10: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Sample/$entry
      -- 
    req_2286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(10), ack => W_tag_1454_delayed_4_0_1524_inst_req_0); -- 
    loadBuffer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(12);
      gj_loadBuffer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: 	24 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Update/req
      -- CP-element group 11: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Update/$entry
      -- CP-element group 11: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_update_start_
      -- 
    req_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(11), ack => W_tag_1454_delayed_4_0_1524_inst_req_1); -- 
    loadBuffer_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(13) & loadBuffer_CP_2250_elements(24);
      gj_loadBuffer_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Sample/ack
      -- CP-element group 12: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Sample/$exit
      -- CP-element group 12: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_sample_completed_
      -- 
    ack_2287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_1454_delayed_4_0_1524_inst_ack_0, ack => loadBuffer_CP_2250_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	22 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Update/ack
      -- CP-element group 13: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_Update/$exit
      -- CP-element group 13: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1526_update_completed_
      -- 
    ack_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_1454_delayed_4_0_1524_inst_ack_1, ack => loadBuffer_CP_2250_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Sample/$entry
      -- CP-element group 14: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Sample/req
      -- CP-element group 14: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_sample_start_
      -- 
    req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(14), ack => W_max_addr_offset_1455_delayed_4_0_1527_inst_req_0); -- 
    loadBuffer_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(16);
      gj_loadBuffer_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	24 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_update_start_
      -- CP-element group 15: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Update/$entry
      -- CP-element group 15: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Update/req
      -- 
    req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(15), ack => W_max_addr_offset_1455_delayed_4_0_1527_inst_req_1); -- 
    loadBuffer_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(17) & loadBuffer_CP_2250_elements(24);
      gj_loadBuffer_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Sample/$exit
      -- CP-element group 16: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Sample/ack
      -- CP-element group 16: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_sample_completed_
      -- 
    ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_max_addr_offset_1455_delayed_4_0_1527_inst_ack_0, ack => loadBuffer_CP_2250_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_update_completed_
      -- CP-element group 17: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Update/$exit
      -- CP-element group 17: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1529_Update/ack
      -- 
    ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_max_addr_offset_1455_delayed_4_0_1527_inst_ack_1, ack => loadBuffer_CP_2250_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: 	9 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_sample_start_
      -- CP-element group 18: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Sample/$entry
      -- CP-element group 18: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Sample/req
      -- 
    req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(18), ack => W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_req_0); -- 
    loadBuffer_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(20);
      gj_loadBuffer_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_update_start_
      -- CP-element group 19: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Update/$entry
      -- CP-element group 19: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Update/req
      -- 
    req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(19), ack => W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_req_1); -- 
    loadBuffer_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(21) & loadBuffer_CP_2250_elements(24);
      gj_loadBuffer_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	4 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_sample_completed_
      -- CP-element group 20: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Sample/ack
      -- 
    ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_ack_0, ack => loadBuffer_CP_2250_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_update_completed_
      -- CP-element group 21: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Update/$exit
      -- CP-element group 21: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1532_Update/ack
      -- 
    ack_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_ack_1, ack => loadBuffer_CP_2250_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	9 
    -- CP-element group 22: 	13 
    -- CP-element group 22: 	17 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_sample_start_
      -- CP-element group 22: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Sample/$entry
      -- CP-element group 22: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Sample/crr
      -- 
    crr_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(22), ack => call_stmt_1540_call_req_0); -- 
    loadBuffer_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(13) & loadBuffer_CP_2250_elements(17) & loadBuffer_CP_2250_elements(21) & loadBuffer_CP_2250_elements(24);
      gj_loadBuffer_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	5 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	44 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_update_start_
      -- CP-element group 23: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Update/ccr
      -- CP-element group 23: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Update/$entry
      -- 
    ccr_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(23), ack => call_stmt_1540_call_req_1); -- 
    loadBuffer_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(5) & loadBuffer_CP_2250_elements(25) & loadBuffer_CP_2250_elements(28) & loadBuffer_CP_2250_elements(44);
      gj_loadBuffer_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	7 
    -- CP-element group 24: 	11 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_sample_completed_
      -- CP-element group 24: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Sample/$exit
      -- CP-element group 24: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Sample/cra
      -- 
    cra_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1540_call_ack_0, ack => loadBuffer_CP_2250_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	42 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_update_completed_
      -- CP-element group 25: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Update/cca
      -- CP-element group 25: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1540_Update/$exit
      -- 
    cca_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1540_call_ack_1, ack => loadBuffer_CP_2250_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	9 
    -- CP-element group 26: 	25 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Sample/req
      -- CP-element group 26: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Sample/$entry
      -- CP-element group 26: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_sample_start_
      -- 
    req_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(26), ack => W_bad_packet_identifier_1462_delayed_8_0_1541_inst_req_0); -- 
    loadBuffer_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(25) & loadBuffer_CP_2250_elements(28);
      gj_loadBuffer_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	44 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Update/req
      -- CP-element group 27: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Update/$entry
      -- CP-element group 27: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_update_start_
      -- 
    req_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(27), ack => W_bad_packet_identifier_1462_delayed_8_0_1541_inst_req_1); -- 
    loadBuffer_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(29) & loadBuffer_CP_2250_elements(44);
      gj_loadBuffer_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Sample/ack
      -- CP-element group 28: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Sample/$exit
      -- CP-element group 28: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_sample_completed_
      -- 
    ack_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1462_delayed_8_0_1541_inst_ack_0, ack => loadBuffer_CP_2250_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	42 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Update/ack
      -- CP-element group 29: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_Update/$exit
      -- CP-element group 29: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1543_update_completed_
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1462_delayed_8_0_1541_inst_ack_1, ack => loadBuffer_CP_2250_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: 	9 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_sample_start_
      -- CP-element group 30: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Sample/$entry
      -- CP-element group 30: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Sample/req
      -- 
    req_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(30), ack => W_tag_1463_delayed_8_0_1544_inst_req_0); -- 
    loadBuffer_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(32);
      gj_loadBuffer_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	44 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_update_start_
      -- CP-element group 31: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Update/$entry
      -- CP-element group 31: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Update/req
      -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(31), ack => W_tag_1463_delayed_8_0_1544_inst_req_1); -- 
    loadBuffer_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(33) & loadBuffer_CP_2250_elements(44);
      gj_loadBuffer_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_sample_completed_
      -- CP-element group 32: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Sample/$exit
      -- CP-element group 32: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Sample/ack
      -- 
    ack_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_1463_delayed_8_0_1544_inst_ack_0, ack => loadBuffer_CP_2250_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	42 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_update_completed_
      -- CP-element group 33: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Update/$exit
      -- CP-element group 33: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1546_Update/ack
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_tag_1463_delayed_8_0_1544_inst_ack_1, ack => loadBuffer_CP_2250_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	1 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_sample_start_
      -- CP-element group 34: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Sample/$entry
      -- CP-element group 34: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Sample/req
      -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(34), ack => W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_req_0); -- 
    loadBuffer_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(36);
      gj_loadBuffer_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	44 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_update_start_
      -- CP-element group 35: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Update/$entry
      -- CP-element group 35: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Update/req
      -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(35), ack => W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_req_1); -- 
    loadBuffer_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(37) & loadBuffer_CP_2250_elements(44);
      gj_loadBuffer_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	4 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_sample_completed_
      -- CP-element group 36: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Sample/$exit
      -- CP-element group 36: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Sample/ack
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_ack_0, ack => loadBuffer_CP_2250_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	42 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_update_completed_
      -- CP-element group 37: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Update/$exit
      -- CP-element group 37: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1549_Update/ack
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_ack_1, ack => loadBuffer_CP_2250_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	1 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_sample_start_
      -- CP-element group 38: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Sample/$entry
      -- CP-element group 38: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Sample/req
      -- 
    req_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(38), ack => W_max_addr_offset_1465_delayed_8_0_1550_inst_req_0); -- 
    loadBuffer_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(1) & loadBuffer_CP_2250_elements(9) & loadBuffer_CP_2250_elements(40);
      gj_loadBuffer_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: 	44 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_update_start_
      -- CP-element group 39: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Update/req
      -- CP-element group 39: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Update/$entry
      -- 
    req_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(39), ack => W_max_addr_offset_1465_delayed_8_0_1550_inst_req_1); -- 
    loadBuffer_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(41) & loadBuffer_CP_2250_elements(44);
      gj_loadBuffer_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	3 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_sample_completed_
      -- CP-element group 40: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Sample/ack
      -- CP-element group 40: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Sample/$exit
      -- 
    ack_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_max_addr_offset_1465_delayed_8_0_1550_inst_ack_0, ack => loadBuffer_CP_2250_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_update_completed_
      -- CP-element group 41: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Update/ack
      -- CP-element group 41: 	 call_stmt_1522_to_call_stmt_1559/assign_stmt_1552_Update/$exit
      -- 
    ack_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_max_addr_offset_1465_delayed_8_0_1550_inst_ack_1, ack => loadBuffer_CP_2250_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	25 
    -- CP-element group 42: 	29 
    -- CP-element group 42: 	33 
    -- CP-element group 42: 	37 
    -- CP-element group 42: 	41 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Sample/crr
      -- CP-element group 42: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Sample/$entry
      -- CP-element group 42: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_sample_start_
      -- 
    crr_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(42), ack => call_stmt_1559_call_req_0); -- 
    loadBuffer_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadBuffer_CP_2250_elements(25) & loadBuffer_CP_2250_elements(29) & loadBuffer_CP_2250_elements(33) & loadBuffer_CP_2250_elements(37) & loadBuffer_CP_2250_elements(41) & loadBuffer_CP_2250_elements(44);
      gj_loadBuffer_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Update/ccr
      -- CP-element group 43: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Update/$entry
      -- CP-element group 43: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_update_start_
      -- 
    ccr_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_2250_elements(43), ack => call_stmt_1559_call_req_1); -- 
    loadBuffer_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_2250_elements(45);
      gj_loadBuffer_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_2250_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	23 
    -- CP-element group 44: 	27 
    -- CP-element group 44: 	31 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	39 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Sample/cra
      -- CP-element group 44: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Sample/$exit
      -- CP-element group 44: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_sample_completed_
      -- 
    cra_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1559_call_ack_0, ack => loadBuffer_CP_2250_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	6 
    -- CP-element group 45: 	43 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Update/cca
      -- CP-element group 45: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_Update/$exit
      -- CP-element group 45: 	 call_stmt_1522_to_call_stmt_1559/call_stmt_1559_update_completed_
      -- CP-element group 45: 	 call_stmt_1522_to_call_stmt_1559/$exit
      -- 
    cca_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1559_call_ack_1, ack => loadBuffer_CP_2250_elements(45)); -- 
    -- CP-element group 46:  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	2 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 tag_update_enable
      -- 
    loadBuffer_CP_2250_elements(46) <= loadBuffer_CP_2250_elements(2);
    -- CP-element group 47:  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	3 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 max_addr_offset_update_enable
      -- 
    loadBuffer_CP_2250_elements(47) <= loadBuffer_CP_2250_elements(3);
    -- CP-element group 48:  place  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	4 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 rx_buffer_pointer_update_enable
      -- 
    loadBuffer_CP_2250_elements(48) <= loadBuffer_CP_2250_elements(4);
    -- CP-element group 49:  place  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	5 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 bad_packet_identifier_update_enable
      -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 $exit
      -- 
    loadBuffer_CP_2250_elements(50) <= loadBuffer_CP_2250_elements(45);
    --  hookup: inputs to control-path 
    loadBuffer_CP_2250_elements(49) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_2250_elements(48);
    max_addr_offset_update_enable <= loadBuffer_CP_2250_elements(47);
    tag_update_enable <= loadBuffer_CP_2250_elements(46);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addr_offset_after_eth_header_1522 : std_logic_vector(15 downto 0);
    signal bad_packet_identifier_1462_delayed_8_0_1543 : std_logic_vector(0 downto 0);
    signal last_keep_1540 : std_logic_vector(7 downto 0);
    signal max_addr_offset_1455_delayed_4_0_1529 : std_logic_vector(15 downto 0);
    signal max_addr_offset_1465_delayed_8_0_1552 : std_logic_vector(15 downto 0);
    signal packet_size_1540 : std_logic_vector(10 downto 0);
    signal rx_buffer_pointer_1456_delayed_4_0_1532 : std_logic_vector(63 downto 0);
    signal rx_buffer_pointer_1464_delayed_8_0_1549 : std_logic_vector(63 downto 0);
    signal tag_1454_delayed_4_0_1526 : std_logic_vector(7 downto 0);
    signal tag_1463_delayed_8_0_1546 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    W_bad_packet_identifier_1462_delayed_8_0_1541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bad_packet_identifier_1462_delayed_8_0_1541_inst_req_0;
      W_bad_packet_identifier_1462_delayed_8_0_1541_inst_ack_0<= wack(0);
      rreq(0) <= W_bad_packet_identifier_1462_delayed_8_0_1541_inst_req_1;
      W_bad_packet_identifier_1462_delayed_8_0_1541_inst_ack_1<= rack(0);
      W_bad_packet_identifier_1462_delayed_8_0_1541_inst : InterlockBuffer generic map ( -- 
        name => "W_bad_packet_identifier_1462_delayed_8_0_1541_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bad_packet_identifier_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bad_packet_identifier_1462_delayed_8_0_1543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_max_addr_offset_1455_delayed_4_0_1527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_max_addr_offset_1455_delayed_4_0_1527_inst_req_0;
      W_max_addr_offset_1455_delayed_4_0_1527_inst_ack_0<= wack(0);
      rreq(0) <= W_max_addr_offset_1455_delayed_4_0_1527_inst_req_1;
      W_max_addr_offset_1455_delayed_4_0_1527_inst_ack_1<= rack(0);
      W_max_addr_offset_1455_delayed_4_0_1527_inst : InterlockBuffer generic map ( -- 
        name => "W_max_addr_offset_1455_delayed_4_0_1527_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => max_addr_offset_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => max_addr_offset_1455_delayed_4_0_1529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_max_addr_offset_1465_delayed_8_0_1550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_max_addr_offset_1465_delayed_8_0_1550_inst_req_0;
      W_max_addr_offset_1465_delayed_8_0_1550_inst_ack_0<= wack(0);
      rreq(0) <= W_max_addr_offset_1465_delayed_8_0_1550_inst_req_1;
      W_max_addr_offset_1465_delayed_8_0_1550_inst_ack_1<= rack(0);
      W_max_addr_offset_1465_delayed_8_0_1550_inst : InterlockBuffer generic map ( -- 
        name => "W_max_addr_offset_1465_delayed_8_0_1550_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => max_addr_offset_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => max_addr_offset_1465_delayed_8_0_1552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_req_0;
      W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_req_1;
      W_rx_buffer_pointer_1456_delayed_4_0_1530_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1456_delayed_4_0_1530_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1456_delayed_4_0_1530_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1456_delayed_4_0_1532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_req_0;
      W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_req_1;
      W_rx_buffer_pointer_1464_delayed_8_0_1547_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1464_delayed_8_0_1547_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1464_delayed_8_0_1547_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1464_delayed_8_0_1549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_tag_1454_delayed_4_0_1524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_tag_1454_delayed_4_0_1524_inst_req_0;
      W_tag_1454_delayed_4_0_1524_inst_ack_0<= wack(0);
      rreq(0) <= W_tag_1454_delayed_4_0_1524_inst_req_1;
      W_tag_1454_delayed_4_0_1524_inst_ack_1<= rack(0);
      W_tag_1454_delayed_4_0_1524_inst : InterlockBuffer generic map ( -- 
        name => "W_tag_1454_delayed_4_0_1524_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_1454_delayed_4_0_1526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_tag_1463_delayed_8_0_1544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_tag_1463_delayed_8_0_1544_inst_req_0;
      W_tag_1463_delayed_8_0_1544_inst_ack_0<= wack(0);
      rreq(0) <= W_tag_1463_delayed_8_0_1544_inst_req_1;
      W_tag_1463_delayed_8_0_1544_inst_ack_1<= rack(0);
      W_tag_1463_delayed_8_0_1544_inst : InterlockBuffer generic map ( -- 
        name => "W_tag_1463_delayed_8_0_1544_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_1463_delayed_8_0_1546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared call operator group (0) : call_stmt_1522_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1522_call_req_0;
      call_stmt_1522_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1522_call_req_1;
      call_stmt_1522_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & rx_buffer_pointer_buffer;
      addr_offset_after_eth_header_1522 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(71 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(15 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1540_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal data_out: std_logic_vector(19 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1540_call_req_0;
      call_stmt_1540_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1540_call_req_1;
      call_stmt_1540_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_1454_delayed_4_0_1526 & max_addr_offset_1455_delayed_4_0_1529 & rx_buffer_pointer_1456_delayed_4_0_1532 & addr_offset_after_eth_header_1522;
      packet_size_1540 <= data_out(19 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_1540 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(103 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 20,
          owidth => 20,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(19 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1559_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(106 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1559_call_req_0;
      call_stmt_1559_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1559_call_req_1;
      call_stmt_1559_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_1462_delayed_8_0_1543(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_1463_delayed_8_0_1546 & rx_buffer_pointer_1464_delayed_8_0_1549 & max_addr_offset_1465_delayed_8_0_1552 & packet_size_1540 & last_keep_1540;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 107,
        owidth => 107,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(106 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_2198_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2206_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_2162_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_2180_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2171_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2177_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2188_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2195_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2204_wire : std_logic_vector(0 downto 0);
    signal MUX_2174_wire : std_logic_vector(1 downto 0);
    signal MUX_2184_wire : std_logic_vector(1 downto 0);
    signal MUX_2191_wire : std_logic_vector(1 downto 0);
    signal MUX_2201_wire : std_logic_vector(1 downto 0);
    signal MUX_2209_wire : std_logic_vector(1 downto 0);
    signal NEQ_u2_u1_2165_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2197_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2181_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_2185_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_2192_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_2210_wire : std_logic_vector(1 downto 0);
    signal R_S0_2170_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_2182_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_2207_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_2172_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_2187_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_2164_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_2189_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_2194_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_2199_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_2203_wire_constant : std_logic_vector(1 downto 0);
    signal R_S3_2176_wire_constant : std_logic_vector(1 downto 0);
    signal go_to_s0_2167 : std_logic_vector(0 downto 0);
    signal konst_2156_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2161_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2173_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2179_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2183_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2190_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2200_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2208_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_2158 : std_logic_vector(0 downto 0);
    signal tlast_2153 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_2170_wire_constant <= "00";
    R_S0_2182_wire_constant <= "00";
    R_S0_2207_wire_constant <= "00";
    R_S1_2172_wire_constant <= "01";
    R_S1_2187_wire_constant <= "01";
    R_S2_2164_wire_constant <= "10";
    R_S2_2189_wire_constant <= "10";
    R_S2_2194_wire_constant <= "10";
    R_S2_2199_wire_constant <= "10";
    R_S2_2203_wire_constant <= "10";
    R_S3_2176_wire_constant <= "11";
    konst_2156_wire_constant <= "1";
    konst_2161_wire_constant <= "1";
    konst_2173_wire_constant <= "00";
    konst_2179_wire_constant <= "1";
    konst_2183_wire_constant <= "00";
    konst_2190_wire_constant <= "00";
    konst_2200_wire_constant <= "00";
    konst_2208_wire_constant <= "00";
    -- flow-through select operator MUX_2174_inst
    MUX_2174_wire <= R_S1_2172_wire_constant when (EQ_u2_u1_2171_wire(0) /=  '0') else konst_2173_wire_constant;
    -- flow-through select operator MUX_2184_inst
    MUX_2184_wire <= R_S0_2182_wire_constant when (OR_u1_u1_2181_wire(0) /=  '0') else konst_2183_wire_constant;
    -- flow-through select operator MUX_2191_inst
    MUX_2191_wire <= R_S2_2189_wire_constant when (EQ_u2_u1_2188_wire(0) /=  '0') else konst_2190_wire_constant;
    -- flow-through select operator MUX_2201_inst
    MUX_2201_wire <= R_S2_2199_wire_constant when (AND_u1_u1_2198_wire(0) /=  '0') else konst_2200_wire_constant;
    -- flow-through select operator MUX_2209_inst
    MUX_2209_wire <= R_S0_2207_wire_constant when (AND_u1_u1_2206_wire(0) /=  '0') else konst_2208_wire_constant;
    -- flow-through slice operator slice_2152_inst
    tlast_2153 <= RX_buffer(72 downto 72);
    -- flow through binary operator AND_u1_u1_2166_inst
    go_to_s0_2167 <= (EQ_u1_u1_2162_wire and NEQ_u2_u1_2165_wire);
    -- flow through binary operator AND_u1_u1_2198_inst
    AND_u1_u1_2198_wire <= (EQ_u2_u1_2195_wire and NOT_u1_u1_2197_wire);
    -- flow through binary operator AND_u1_u1_2206_inst
    AND_u1_u1_2206_wire <= (EQ_u2_u1_2204_wire and last_word_2158);
    -- flow through binary operator EQ_u1_u1_2157_inst
    process(tlast_2153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_2153, konst_2156_wire_constant, tmp_var);
      last_word_2158 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_2162_inst
    process(last_word_2158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_word_2158, konst_2161_wire_constant, tmp_var);
      EQ_u1_u1_2162_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u1_u1_2180_inst
    process(go_to_s0_2167) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(go_to_s0_2167, konst_2179_wire_constant, tmp_var);
      EQ_u1_u1_2180_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2171_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_2170_wire_constant, tmp_var);
      EQ_u2_u1_2171_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2177_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S3_2176_wire_constant, tmp_var);
      EQ_u2_u1_2177_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2188_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_2187_wire_constant, tmp_var);
      EQ_u2_u1_2188_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2195_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_2194_wire_constant, tmp_var);
      EQ_u2_u1_2195_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2204_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_2203_wire_constant, tmp_var);
      EQ_u2_u1_2204_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u2_u1_2165_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSTATE_buffer, R_S2_2164_wire_constant, tmp_var);
      NEQ_u2_u1_2165_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2197_inst
    process(last_word_2158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_2158, tmp_var);
      NOT_u1_u1_2197_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_2181_inst
    OR_u1_u1_2181_wire <= (EQ_u2_u1_2177_wire or EQ_u1_u1_2180_wire);
    -- flow through binary operator OR_u2_u2_2185_inst
    OR_u2_u2_2185_wire <= (MUX_2174_wire or MUX_2184_wire);
    -- flow through binary operator OR_u2_u2_2192_inst
    OR_u2_u2_2192_wire <= (OR_u2_u2_2185_wire or MUX_2191_wire);
    -- flow through binary operator OR_u2_u2_2210_inst
    OR_u2_u2_2210_wire <= (MUX_2201_wire or MUX_2209_wire);
    -- flow through binary operator OR_u2_u2_2211_inst
    nLSTATE_buffer <= (OR_u2_u2_2192_wire or OR_u2_u2_2210_wire);
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    S_CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(1 downto 0);
    accessRegister_call_acks : in   std_logic_vector(1 downto 0);
    accessRegister_call_data : out  std_logic_vector(89 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(1 downto 0);
    accessRegister_return_acks : in   std_logic_vector(1 downto 0);
    accessRegister_return_data : in   std_logic_vector(63 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_4047_start: Boolean;
  signal nicRxFromMacDaemon_CP_4047_symbol: Boolean;
  -- volatile/operator module components. 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component nextLSTATE_Volatile is -- 
    port ( -- 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal if_stmt_2228_branch_ack_0 : boolean;
  signal npkt_cnt_2305_2259_buf_req_1 : boolean;
  signal call_stmt_2245_call_req_1 : boolean;
  signal call_stmt_2245_call_ack_1 : boolean;
  signal nLSTATE_2267_2250_buf_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_2254_inst_ack_0 : boolean;
  signal nLSTATE_2267_2250_buf_req_1 : boolean;
  signal if_stmt_2228_branch_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_2254_inst_ack_1 : boolean;
  signal call_stmt_2245_call_ack_0 : boolean;
  signal phi_stmt_2248_ack_0 : boolean;
  signal nLSTATE_2267_2250_buf_ack_1 : boolean;
  signal call_stmt_2245_call_req_0 : boolean;
  signal phi_stmt_2255_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_2254_inst_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_2254_inst_req_0 : boolean;
  signal phi_stmt_2248_req_0 : boolean;
  signal do_while_stmt_2246_branch_req_0 : boolean;
  signal if_stmt_2228_branch_ack_1 : boolean;
  signal MUX_2287_inst_ack_1 : boolean;
  signal phi_stmt_2255_req_1 : boolean;
  signal npkt_cnt_2305_2259_buf_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_2278_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_2278_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_2289_inst_req_0 : boolean;
  signal call_stmt_2315_call_req_1 : boolean;
  signal WPIPE_nic_rx_to_packet_2289_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_packet_2289_inst_ack_1 : boolean;
  signal call_stmt_2315_call_ack_1 : boolean;
  signal MUX_2287_inst_ack_0 : boolean;
  signal MUX_2287_inst_req_0 : boolean;
  signal npkt_cnt_2305_2259_buf_ack_0 : boolean;
  signal npkt_cnt_2305_2259_buf_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_2278_inst_req_1 : boolean;
  signal MUX_2287_inst_req_1 : boolean;
  signal phi_stmt_2248_req_1 : boolean;
  signal phi_stmt_2255_req_0 : boolean;
  signal do_while_stmt_2246_branch_ack_0 : boolean;
  signal do_while_stmt_2246_branch_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_2278_inst_ack_1 : boolean;
  signal call_stmt_2315_call_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_2289_inst_ack_0 : boolean;
  signal call_stmt_2315_call_req_0 : boolean;
  signal nLSTATE_2267_2250_buf_ack_0 : boolean;
  signal call_stmt_2227_call_req_0 : boolean;
  signal call_stmt_2227_call_ack_0 : boolean;
  signal call_stmt_2227_call_req_1 : boolean;
  signal call_stmt_2227_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_4047_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_4047_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_4047_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_4047_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_4047: Block -- control-path 
    signal nicRxFromMacDaemon_CP_4047_elements: BooleanArray(83 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_4047_elements(0) <= nicRxFromMacDaemon_CP_4047_start;
    nicRxFromMacDaemon_CP_4047_symbol <= nicRxFromMacDaemon_CP_4047_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	83 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_2215/merge_stmt_2217__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/merge_stmt_2217__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_2215/merge_stmt_2217_dead_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2215/$entry
      -- CP-element group 0: 	 branch_block_stmt_2215/branch_block_stmt_2215__entry__
      -- CP-element group 0: 	 branch_block_stmt_2215/merge_stmt_2217__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2215/$exit
      -- CP-element group 1: 	 branch_block_stmt_2215/branch_block_stmt_2215__exit__
      -- 
    nicRxFromMacDaemon_CP_4047_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	82 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	83 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_2215/disable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_2215/disable_loopback_PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_2215/do_while_stmt_2246__exit__
      -- CP-element group 2: 	 branch_block_stmt_2215/disable_loopback
      -- 
    nicRxFromMacDaemon_CP_4047_elements(2) <= nicRxFromMacDaemon_CP_4047_elements(82);
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	83 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Sample/cra
      -- 
    cra_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2227_call_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	83 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (49) 
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_else_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2215/NOT_u1_u1_2232_place
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/call_stmt_2227__exit__
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228__entry__
      -- CP-element group 4: 	 branch_block_stmt_2215/call_stmt_2227/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Sample/req
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Sample/ack
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Update/req
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/BITSEL_u32_u1_2231_inputs/RPIPE_S_CONTROL_REGISTER_2229/Update/ack
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/BITSEL_u32_u1_2231/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2215/if_stmt_2228_eval_test/NOT_u1_u1_2232/SplitProtocol/Update/$entry
      -- 
    cca_4082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2227_call_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(4)); -- 
    branch_req_4138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(4), ack => if_stmt_2228_branch_req_0); -- 
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	83 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2215/if_stmt_2228_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_2215/if_stmt_2228_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_2215/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_2215/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_2215/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_4143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2228_branch_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(5)); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_2215/if_stmt_2228_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_2215/if_stmt_2228_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Update/ccr
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/$entry
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2215/if_stmt_2228__exit__
      -- CP-element group 6: 	 branch_block_stmt_2215/call_stmt_2245__entry__
      -- 
    else_choice_transition_4147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2228_branch_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(6)); -- 
    ccr_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(6), ack => call_stmt_2245_call_req_1); -- 
    crr_4159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(6), ack => call_stmt_2245_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Sample/cra
      -- CP-element group 7: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_sample_completed_
      -- 
    cra_4160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2245_call_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Update/cca
      -- CP-element group 8: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2215/call_stmt_2245/$exit
      -- CP-element group 8: 	 branch_block_stmt_2215/call_stmt_2245/call_stmt_2245_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2215/call_stmt_2245__exit__
      -- CP-element group 8: 	 branch_block_stmt_2215/do_while_stmt_2246__entry__
      -- 
    cca_4165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2245_call_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(8)); -- 
    -- CP-element group 9:  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246__entry__
      -- CP-element group 9: 	 branch_block_stmt_2215/do_while_stmt_2246/$entry
      -- 
    nicRxFromMacDaemon_CP_4047_elements(9) <= nicRxFromMacDaemon_CP_4047_elements(8);
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	82 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246__exit__
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(10) is bound as output of CP function.
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_back
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(11) is bound as output of CP function.
    -- CP-element group 12:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	80 
    -- CP-element group 12: 	81 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2215/do_while_stmt_2246/condition_done
      -- CP-element group 12: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_exit/$entry
      -- CP-element group 12: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_taken/$entry
      -- 
    nicRxFromMacDaemon_CP_4047_elements(12) <= nicRxFromMacDaemon_CP_4047_elements(17);
    -- CP-element group 13:  branch  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	79 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_body_done
      -- 
    nicRxFromMacDaemon_CP_4047_elements(13) <= nicRxFromMacDaemon_CP_4047_elements(79);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14: 	51 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/back_edge_to_loop_body
      -- 
    nicRxFromMacDaemon_CP_4047_elements(14) <= nicRxFromMacDaemon_CP_4047_elements(11);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	53 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/first_time_through_loop_body
      -- 
    nicRxFromMacDaemon_CP_4047_elements(15) <= nicRxFromMacDaemon_CP_4047_elements(9);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	23 
    -- CP-element group 16: 	24 
    -- CP-element group 16: 	40 
    -- CP-element group 16: 	45 
    -- CP-element group 16: 	46 
    -- CP-element group 16: 	78 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/loop_body_start
      -- CP-element group 16: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2252_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/$entry
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(16) is bound as output of CP function.
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	78 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/condition_evaluated
      -- 
    condition_evaluated_4180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(17), ack => do_while_stmt_2246_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(22) & nicRxFromMacDaemon_CP_4047_elements(78);
      gj_nicRxFromMacDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	45 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	47 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_sample_start__ps
      -- CP-element group 18: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/aggregated_phi_sample_req
      -- 
    nicRxFromMacDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(16) & nicRxFromMacDaemon_CP_4047_elements(23) & nicRxFromMacDaemon_CP_4047_elements(45) & nicRxFromMacDaemon_CP_4047_elements(22);
      gj_nicRxFromMacDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	25 
    -- CP-element group 19: 	43 
    -- CP-element group 19: 	48 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	79 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	45 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2252_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_sample_completed_
      -- 
    nicRxFromMacDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(25) & nicRxFromMacDaemon_CP_4047_elements(43) & nicRxFromMacDaemon_CP_4047_elements(48);
      gj_nicRxFromMacDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	79 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(20) is a control-delay.
    cp_element_20_delay: control_delay_element  generic map(name => " 20_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_4047_elements(19), ack => nicRxFromMacDaemon_CP_4047_elements(20), clk => clk, reset =>reset);
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	40 
    -- CP-element group 21: 	46 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	42 
    -- CP-element group 21: 	49 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_update_start__ps
      -- CP-element group 21: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/aggregated_phi_update_req
      -- 
    nicRxFromMacDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(24) & nicRxFromMacDaemon_CP_4047_elements(40) & nicRxFromMacDaemon_CP_4047_elements(46);
      gj_nicRxFromMacDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: 	44 
    -- CP-element group 22: 	50 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/aggregated_phi_update_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(26) & nicRxFromMacDaemon_CP_4047_elements(44) & nicRxFromMacDaemon_CP_4047_elements(50);
      gj_nicRxFromMacDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	18 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(16) & nicRxFromMacDaemon_CP_4047_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	16 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	66 
    -- CP-element group 24: 	69 
    -- CP-element group 24: 	76 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	21 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(16) & nicRxFromMacDaemon_CP_4047_elements(26) & nicRxFromMacDaemon_CP_4047_elements(66) & nicRxFromMacDaemon_CP_4047_elements(69) & nicRxFromMacDaemon_CP_4047_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	19 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: 	64 
    -- CP-element group 26: 	68 
    -- CP-element group 26: 	74 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_update_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_4047_elements(27) <= nicRxFromMacDaemon_CP_4047_elements(14);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_loopback_sample_req
      -- CP-element group 28: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_loopback_sample_req_ps
      -- 
    phi_stmt_2248_loopback_sample_req_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2248_loopback_sample_req_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(28), ack => phi_stmt_2248_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_4047_elements(29) <= nicRxFromMacDaemon_CP_4047_elements(15);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_entry_sample_req_ps
      -- CP-element group 30: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_entry_sample_req
      -- 
    phi_stmt_2248_entry_sample_req_4199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2248_entry_sample_req_4199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(30), ack => phi_stmt_2248_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_phi_mux_ack
      -- CP-element group 31: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2248_phi_mux_ack_ps
      -- 
    phi_stmt_2248_phi_mux_ack_4202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2248_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Sample/req
      -- CP-element group 32: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_sample_start__ps
      -- 
    req_4215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(32), ack => nLSTATE_2267_2250_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Update/req
      -- CP-element group 33: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_update_start_
      -- CP-element group 33: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_update_start__ps
      -- 
    req_4220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(33), ack => nLSTATE_2267_2250_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Sample/ack
      -- 
    ack_4216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_2267_2250_buf_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_nLSTATE_2250_Update/ack
      -- 
    ack_4221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_2267_2250_buf_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_sample_start__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_update_start_
      -- CP-element group 37: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_update_start__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_4047_elements(38) <= nicRxFromMacDaemon_CP_4047_elements(39);
    -- CP-element group 39:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	38 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_S0_2251_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(39) is a control-delay.
    cp_element_39_delay: control_delay_element  generic map(name => " 39_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_4047_elements(37), ack => nicRxFromMacDaemon_CP_4047_elements(39), clk => clk, reset =>reset);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	16 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	66 
    -- CP-element group 40: 	72 
    -- CP-element group 40: 	76 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	21 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2252_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(16) & nicRxFromMacDaemon_CP_4047_elements(66) & nicRxFromMacDaemon_CP_4047_elements(72) & nicRxFromMacDaemon_CP_4047_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	44 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Sample/$entry
      -- 
    rr_4242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(41), ack => RPIPE_mac_to_nic_data_2254_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(18) & nicRxFromMacDaemon_CP_4047_elements(44);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	21 
    -- CP-element group 42: 	43 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_update_start_
      -- CP-element group 42: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Update/cr
      -- 
    cr_4247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(42), ack => RPIPE_mac_to_nic_data_2254_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(21) & nicRxFromMacDaemon_CP_4047_elements(43);
      gj_nicRxFromMacDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	19 
    -- CP-element group 43: 	42 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Sample/$exit
      -- 
    ra_4243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_2254_inst_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	22 
    -- CP-element group 44: 	64 
    -- CP-element group 44: 	71 
    -- CP-element group 44: 	74 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	41 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2252_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/RPIPE_mac_to_nic_data_2254_Update/$exit
      -- 
    ca_4248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_2254_inst_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(44)); -- 
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	16 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	19 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	18 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(16) & nicRxFromMacDaemon_CP_4047_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	50 
    -- CP-element group 46: 	76 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	21 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(16) & nicRxFromMacDaemon_CP_4047_elements(50) & nicRxFromMacDaemon_CP_4047_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	18 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_sample_start__ps
      -- 
    nicRxFromMacDaemon_CP_4047_elements(47) <= nicRxFromMacDaemon_CP_4047_elements(18);
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	19 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	21 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_update_start__ps
      -- 
    nicRxFromMacDaemon_CP_4047_elements(49) <= nicRxFromMacDaemon_CP_4047_elements(21);
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	22 
    -- CP-element group 50: 	74 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	46 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(50) is bound as output of CP function.
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	14 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_4047_elements(51) <= nicRxFromMacDaemon_CP_4047_elements(14);
    -- CP-element group 52:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_loopback_sample_req
      -- CP-element group 52: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_loopback_sample_req_ps
      -- 
    phi_stmt_2255_loopback_sample_req_4258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2255_loopback_sample_req_4258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(52), ack => phi_stmt_2255_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(52) is bound as output of CP function.
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	15 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_4047_elements(53) <= nicRxFromMacDaemon_CP_4047_elements(15);
    -- CP-element group 54:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_entry_sample_req_ps
      -- CP-element group 54: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_entry_sample_req
      -- 
    phi_stmt_2255_entry_sample_req_4261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2255_entry_sample_req_4261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(54), ack => phi_stmt_2255_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_phi_mux_ack_ps
      -- CP-element group 55: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/phi_stmt_2255_phi_mux_ack
      -- 
    phi_stmt_2255_phi_mux_ack_4264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2255_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_sample_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_sample_start__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_4047_elements(58) <= nicRxFromMacDaemon_CP_4047_elements(59);
    -- CP-element group 59:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	58 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/type_cast_2258_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(59) is a control-delay.
    cp_element_59_delay: control_delay_element  generic map(name => " 59_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_4047_elements(57), ack => nicRxFromMacDaemon_CP_4047_elements(59), clk => clk, reset =>reset);
    -- CP-element group 60:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (4) 
      -- CP-element group 60: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_sample_start__ps
      -- 
    req_4285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(60), ack => npkt_cnt_2305_2259_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Update/req
      -- CP-element group 61: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_update_start_
      -- CP-element group 61: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_update_start__ps
      -- 
    req_4290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(61), ack => npkt_cnt_2305_2259_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Sample/ack
      -- CP-element group 62: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_sample_completed__ps
      -- 
    ack_4286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_2305_2259_buf_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(62)); -- 
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_Update/ack
      -- CP-element group 63: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/R_npkt_cnt_2259_update_completed__ps
      -- 
    ack_4291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_2305_2259_buf_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	26 
    -- CP-element group 64: 	44 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_start/req
      -- CP-element group 64: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_sample_start_
      -- 
    req_4300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(64), ack => MUX_2287_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(26) & nicRxFromMacDaemon_CP_4047_elements(44) & nicRxFromMacDaemon_CP_4047_elements(66);
      gj_nicRxFromMacDaemon_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	69 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_complete/req
      -- 
    req_4305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(65), ack => MUX_2287_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(67) & nicRxFromMacDaemon_CP_4047_elements(69);
      gj_nicRxFromMacDaemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	24 
    -- CP-element group 66: 	40 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_start/ack
      -- CP-element group 66: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_start/$exit
      -- CP-element group 66: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_sample_completed_
      -- 
    ack_4301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2287_inst_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_complete/ack
      -- CP-element group 67: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/MUX_2287_complete/$exit
      -- 
    ack_4306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2287_inst_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	26 
    -- CP-element group 68: 	67 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Sample/req
      -- CP-element group 68: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_sample_start_
      -- 
    req_4314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(68), ack => WPIPE_nic_rx_to_header_2278_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(26) & nicRxFromMacDaemon_CP_4047_elements(67) & nicRxFromMacDaemon_CP_4047_elements(70);
      gj_nicRxFromMacDaemon_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	24 
    -- CP-element group 69: 	65 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Update/req
      -- CP-element group 69: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Update/$entry
      -- 
    ack_4315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_2278_inst_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(69)); -- 
    req_4319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(69), ack => WPIPE_nic_rx_to_header_2278_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	79 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_header_2278_Update/ack
      -- 
    ack_4320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_2278_inst_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	44 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_sample_start_
      -- 
    req_4328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(71), ack => WPIPE_nic_rx_to_packet_2289_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(44) & nicRxFromMacDaemon_CP_4047_elements(73);
      gj_nicRxFromMacDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	40 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_update_start_
      -- CP-element group 72: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Update/req
      -- CP-element group 72: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Sample/ack
      -- 
    ack_4329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_2289_inst_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(72)); -- 
    req_4333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(72), ack => WPIPE_nic_rx_to_packet_2289_inst_req_1); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	79 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/WPIPE_nic_rx_to_packet_2289_Update/$exit
      -- 
    ack_4334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_2289_inst_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	26 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	50 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Sample/crr
      -- 
    crr_4342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(74), ack => call_stmt_2315_call_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(26) & nicRxFromMacDaemon_CP_4047_elements(44) & nicRxFromMacDaemon_CP_4047_elements(50) & nicRxFromMacDaemon_CP_4047_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Update/ccr
      -- CP-element group 75: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Update/$entry
      -- 
    ccr_4347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(75), ack => call_stmt_2315_call_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicRxFromMacDaemon_CP_4047_elements(77);
      gj_nicRxFromMacDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	24 
    -- CP-element group 76: 	40 
    -- CP-element group 76: 	46 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Sample/cra
      -- CP-element group 76: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Sample/$exit
      -- 
    cra_4343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2315_call_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_Update/cca
      -- CP-element group 77: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/call_stmt_2315_update_completed_
      -- 
    cca_4348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2315_call_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(77)); -- 
    -- CP-element group 78:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	16 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	17 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_4047_elements(78) is a control-delay.
    cp_element_78_delay: control_delay_element  generic map(name => " 78_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_4047_elements(16), ack => nicRxFromMacDaemon_CP_4047_elements(78), clk => clk, reset =>reset);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	19 
    -- CP-element group 79: 	20 
    -- CP-element group 79: 	70 
    -- CP-element group 79: 	73 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	13 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2215/do_while_stmt_2246/do_while_stmt_2246_loop_body/$exit
      -- 
    nicRxFromMacDaemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_4047_elements(19) & nicRxFromMacDaemon_CP_4047_elements(20) & nicRxFromMacDaemon_CP_4047_elements(70) & nicRxFromMacDaemon_CP_4047_elements(73) & nicRxFromMacDaemon_CP_4047_elements(77);
      gj_nicRxFromMacDaemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	12 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_exit/$exit
      -- CP-element group 80: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_exit/ack
      -- 
    ack_4353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2246_branch_ack_0, ack => nicRxFromMacDaemon_CP_4047_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	12 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_taken/$exit
      -- CP-element group 81: 	 branch_block_stmt_2215/do_while_stmt_2246/loop_taken/ack
      -- 
    ack_4357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2246_branch_ack_1, ack => nicRxFromMacDaemon_CP_4047_elements(81)); -- 
    -- CP-element group 82:  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	10 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	2 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2215/do_while_stmt_2246/$exit
      -- 
    nicRxFromMacDaemon_CP_4047_elements(82) <= nicRxFromMacDaemon_CP_4047_elements(10);
    -- CP-element group 83:  merge  fork  transition  place  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	0 
    -- CP-element group 83: 	2 
    -- CP-element group 83: 	5 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	3 
    -- CP-element group 83: 	4 
    -- CP-element group 83:  members (13) 
      -- CP-element group 83: 	 branch_block_stmt_2215/merge_stmt_2217_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_2215/merge_stmt_2217_PhiAck/$entry
      -- CP-element group 83: 	 branch_block_stmt_2215/merge_stmt_2217_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_2215/merge_stmt_2217__exit__
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227__entry__
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/$entry
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_update_start_
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Sample/crr
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_2215/call_stmt_2227/call_stmt_2227_Update/ccr
      -- CP-element group 83: 	 branch_block_stmt_2215/merge_stmt_2217_PhiAck/dummy
      -- 
    crr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(83), ack => call_stmt_2227_call_req_0); -- 
    ccr_4081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_4047_elements(83), ack => call_stmt_2227_call_req_1); -- 
    nicRxFromMacDaemon_CP_4047_elements(83) <= OrReduce(nicRxFromMacDaemon_CP_4047_elements(0) & nicRxFromMacDaemon_CP_4047_elements(2) & nicRxFromMacDaemon_CP_4047_elements(5));
    nicRxFromMacDaemon_do_while_stmt_2246_terminator_4358: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_2246_terminator_4358", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_4047_elements(13),loop_continue => nicRxFromMacDaemon_CP_4047_elements(81),loop_terminate => nicRxFromMacDaemon_CP_4047_elements(80),loop_back => nicRxFromMacDaemon_CP_4047_elements(11),loop_exit => nicRxFromMacDaemon_CP_4047_elements(10),clk => clk, reset => reset); -- 
    phi_stmt_2248_phi_seq_4230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_4047_elements(27);
      nicRxFromMacDaemon_CP_4047_elements(32)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_4047_elements(34);
      nicRxFromMacDaemon_CP_4047_elements(33)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_4047_elements(35);
      nicRxFromMacDaemon_CP_4047_elements(28) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_4047_elements(29);
      nicRxFromMacDaemon_CP_4047_elements(36)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_4047_elements(36);
      nicRxFromMacDaemon_CP_4047_elements(37)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_4047_elements(38);
      nicRxFromMacDaemon_CP_4047_elements(30) <= phi_mux_reqs(1);
      phi_stmt_2248_phi_seq_4230 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2248_phi_seq_4230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_4047_elements(18), 
          phi_sample_ack => nicRxFromMacDaemon_CP_4047_elements(25), 
          phi_update_req => nicRxFromMacDaemon_CP_4047_elements(21), 
          phi_update_ack => nicRxFromMacDaemon_CP_4047_elements(26), 
          phi_mux_ack => nicRxFromMacDaemon_CP_4047_elements(31), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2255_phi_seq_4292_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_4047_elements(53);
      nicRxFromMacDaemon_CP_4047_elements(56)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_4047_elements(56);
      nicRxFromMacDaemon_CP_4047_elements(57)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_4047_elements(58);
      nicRxFromMacDaemon_CP_4047_elements(54) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_4047_elements(51);
      nicRxFromMacDaemon_CP_4047_elements(60)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_4047_elements(62);
      nicRxFromMacDaemon_CP_4047_elements(61)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_4047_elements(63);
      nicRxFromMacDaemon_CP_4047_elements(52) <= phi_mux_reqs(1);
      phi_stmt_2255_phi_seq_4292 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2255_phi_seq_4292") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_4047_elements(47), 
          phi_sample_ack => nicRxFromMacDaemon_CP_4047_elements(48), 
          phi_update_req => nicRxFromMacDaemon_CP_4047_elements(49), 
          phi_update_ack => nicRxFromMacDaemon_CP_4047_elements(50), 
          phi_mux_ack => nicRxFromMacDaemon_CP_4047_elements(55), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4181_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_4047_elements(14);
        preds(1)  <= nicRxFromMacDaemon_CP_4047_elements(15);
        entry_tmerge_4181 : transition_merge -- 
          generic map(name => " entry_tmerge_4181")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_4047_elements(16));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_2302_wire : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_2231_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2322_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u65_u73_2285_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_2271_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2274_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2281_wire : std_logic_vector(0 downto 0);
    signal LSTATE_2248 : std_logic_vector(1 downto 0);
    signal MUX_2287_wire : std_logic_vector(72 downto 0);
    signal NOT_u1_u1_2232_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_2222_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_2240_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_2311_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_S_CONTROL_REGISTER_2229_wire : std_logic_vector(31 downto 0);
    signal RPIPE_S_CONTROL_REGISTER_2320_wire : std_logic_vector(31 downto 0);
    signal RPIPE_mac_to_nic_data_2254_wire : std_logic_vector(72 downto 0);
    signal RX_2252 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_2284_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_2251_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_2270_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_2294_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_2273_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_2280_wire_constant : std_logic_vector(1 downto 0);
    signal ignore_resp0_2227 : std_logic_vector(31 downto 0);
    signal ignore_resp1_2245 : std_logic_vector(31 downto 0);
    signal ignore_resp2_2315 : std_logic_vector(31 downto 0);
    signal konst_2223_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2230_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2241_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2312_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2321_wire_constant : std_logic_vector(31 downto 0);
    signal nLSTATE_2267 : std_logic_vector(1 downto 0);
    signal nLSTATE_2267_2250_buffered : std_logic_vector(1 downto 0);
    signal npkt_cnt_2305 : std_logic_vector(31 downto 0);
    signal npkt_cnt_2305_2259_buffered : std_logic_vector(31 downto 0);
    signal pkt_cnt_2255 : std_logic_vector(31 downto 0);
    signal pkt_complete_2296 : std_logic_vector(0 downto 0);
    signal slice_2283_wire : std_logic_vector(64 downto 0);
    signal type_cast_2219_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2225_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2237_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2243_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2258_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2301_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2308_wire_constant : std_logic_vector(0 downto 0);
    signal write_to_header_2276 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_2222_wire_constant <= "1111";
    NOT_u4_u4_2240_wire_constant <= "1111";
    NOT_u4_u4_2311_wire_constant <= "1111";
    R_HEADER_TKEEP_2284_wire_constant <= "11111100";
    R_S0_2251_wire_constant <= "00";
    R_S0_2270_wire_constant <= "00";
    R_S0_2294_wire_constant <= "00";
    R_S1_2273_wire_constant <= "01";
    R_S1_2280_wire_constant <= "01";
    konst_2223_wire_constant <= "00010110";
    konst_2230_wire_constant <= "00000000000000000000000000000000";
    konst_2241_wire_constant <= "11010100";
    konst_2312_wire_constant <= "00010111";
    konst_2321_wire_constant <= "00000000000000000000000000000000";
    type_cast_2219_wire_constant <= "0";
    type_cast_2225_wire_constant <= "00000000000000000000000000000000";
    type_cast_2237_wire_constant <= "0";
    type_cast_2243_wire_constant <= "00000000000000000000000000000001";
    type_cast_2258_wire_constant <= "00000000000000000000000000000000";
    type_cast_2301_wire_constant <= "00000000000000000000000000000001";
    type_cast_2308_wire_constant <= "0";
    phi_stmt_2248: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nLSTATE_2267_2250_buffered & R_S0_2251_wire_constant;
      req <= phi_stmt_2248_req_0 & phi_stmt_2248_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2248",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2248_ack_0,
          idata => idata,
          odata => LSTATE_2248,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2248
    phi_stmt_2255: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2258_wire_constant & npkt_cnt_2305_2259_buffered;
      req <= phi_stmt_2255_req_0 & phi_stmt_2255_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2255",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2255_ack_0,
          idata => idata,
          odata => pkt_cnt_2255,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2255
    MUX_2287_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_2287_inst_req_0;
      MUX_2287_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_2287_inst_req_1;
      MUX_2287_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_2276(0);
      MUX_2287_inst_gI: SplitGuardInterface generic map(name => "MUX_2287_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_2287_inst: SelectSplitProtocol generic map(name => "MUX_2287_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_2285_wire, y => RX_2252, sel => EQ_u2_u1_2281_wire, z => MUX_2287_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_2304_inst
    npkt_cnt_2305 <= ADD_u32_u32_2302_wire when (pkt_complete_2296(0) /=  '0') else pkt_cnt_2255;
    -- flow-through slice operator slice_2283_inst
    slice_2283_wire <= RX_2252(72 downto 8);
    nLSTATE_2267_2250_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_2267_2250_buf_req_0;
      nLSTATE_2267_2250_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_2267_2250_buf_req_1;
      nLSTATE_2267_2250_buf_ack_1<= rack(0);
      nLSTATE_2267_2250_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_2267_2250_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_2267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_2267_2250_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_2305_2259_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_2305_2259_buf_req_0;
      npkt_cnt_2305_2259_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_2305_2259_buf_req_1;
      npkt_cnt_2305_2259_buf_ack_1<= rack(0);
      npkt_cnt_2305_2259_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_2305_2259_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_2305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_2305_2259_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2252
    process(RPIPE_mac_to_nic_data_2254_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_2254_wire(72 downto 0);
      RX_2252 <= tmp_var; -- 
    end process;
    do_while_stmt_2246_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_2322_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2246_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2246_branch_req_0,
          ack0 => do_while_stmt_2246_branch_ack_0,
          ack1 => do_while_stmt_2246_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2228_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2232_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2228_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2228_branch_req_0,
          ack0 => if_stmt_2228_branch_ack_0,
          ack1 => if_stmt_2228_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u32_u32_2302_inst
    ADD_u32_u32_2302_wire <= std_logic_vector(unsigned(pkt_cnt_2255) + unsigned(type_cast_2301_wire_constant));
    -- flow through binary operator BITSEL_u32_u1_2231_inst
    process(RPIPE_S_CONTROL_REGISTER_2229_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_S_CONTROL_REGISTER_2229_wire, konst_2230_wire_constant, tmp_var);
      BITSEL_u32_u1_2231_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_2322_inst
    process(RPIPE_S_CONTROL_REGISTER_2320_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_S_CONTROL_REGISTER_2320_wire, konst_2321_wire_constant, tmp_var);
      BITSEL_u32_u1_2322_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u65_u73_2285_inst
    process(slice_2283_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_2283_wire, R_HEADER_TKEEP_2284_wire_constant, tmp_var);
      CONCAT_u65_u73_2285_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2271_inst
    process(LSTATE_2248) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_2248, R_S0_2270_wire_constant, tmp_var);
      EQ_u2_u1_2271_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2274_inst
    process(LSTATE_2248) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_2248, R_S1_2273_wire_constant, tmp_var);
      EQ_u2_u1_2274_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2281_inst
    process(LSTATE_2248) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_2248, R_S1_2280_wire_constant, tmp_var);
      EQ_u2_u1_2281_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u2_u1_2295_inst
    process(nLSTATE_2267) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(nLSTATE_2267, R_S0_2294_wire_constant, tmp_var);
      pkt_complete_2296 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2232_inst
    process(BITSEL_u32_u1_2231_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_2231_wire, tmp_var);
      NOT_u1_u1_2232_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_2275_inst
    write_to_header_2276 <= (EQ_u2_u1_2271_wire or EQ_u2_u1_2274_wire);
    -- read from input-signal S_CONTROL_REGISTER
    RPIPE_S_CONTROL_REGISTER_2229_wire <= S_CONTROL_REGISTER;
    -- read from input-signal S_CONTROL_REGISTER
    RPIPE_S_CONTROL_REGISTER_2320_wire <= S_CONTROL_REGISTER;
    -- shared inport operator group (2) : RPIPE_mac_to_nic_data_2254_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_2254_inst_req_0;
      RPIPE_mac_to_nic_data_2254_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_2254_inst_req_1;
      RPIPE_mac_to_nic_data_2254_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_2254_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_2_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_2: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_2", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_2278_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_2278_inst_req_0;
      WPIPE_nic_rx_to_header_2278_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_2278_inst_req_1;
      WPIPE_nic_rx_to_header_2278_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_2276(0);
      data_in <= MUX_2287_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_2289_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_2289_inst_req_0;
      WPIPE_nic_rx_to_packet_2289_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_2289_inst_req_1;
      WPIPE_nic_rx_to_packet_2289_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_2252;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2227_call call_stmt_2245_call 
    accessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2227_call_req_0;
      reqL_unguarded(0) <= call_stmt_2245_call_req_0;
      call_stmt_2227_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2245_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2227_call_req_1;
      reqR_unguarded(0) <= call_stmt_2245_call_req_1;
      call_stmt_2227_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2245_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2219_wire_constant & NOT_u4_u4_2222_wire_constant & konst_2223_wire_constant & type_cast_2225_wire_constant & type_cast_2237_wire_constant & NOT_u4_u4_2240_wire_constant & konst_2241_wire_constant & type_cast_2243_wire_constant;
      ignore_resp0_2227 <= data_out(63 downto 32);
      ignore_resp1_2245 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 90,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(1),
          ackR => accessRegister_call_acks(1),
          dataR => accessRegister_call_data(89 downto 45),
          tagR => accessRegister_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(1), -- cross-over
          ackL => accessRegister_return_reqs(1), -- cross-over
          dataL => accessRegister_return_data(63 downto 32),
          tagL => accessRegister_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_nextLSTATE_6265: nextLSTATE_Volatile port map(RX => RX_2252, LSTATE => LSTATE_2248, nLSTATE => nLSTATE_2267); 
    -- shared call operator group (2) : call_stmt_2315_call 
    accessRegister_call_group_2: Block -- 
      signal data_in: std_logic_vector(44 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2315_call_req_0;
      call_stmt_2315_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2315_call_req_1;
      call_stmt_2315_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= pkt_complete_2296(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessRegister_call_group_2_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2308_wire_constant & NOT_u4_u4_2311_wire_constant & konst_2312_wire_constant & pkt_cnt_2255;
      ignore_resp2_2315 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 45,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    queue_type : in  std_logic_vector(1 downto 0);
    server_id : in  std_logic_vector(7 downto 0);
    q_r_data : out  std_logic_vector(63 downto 0);
    status : out  std_logic_vector(0 downto 0);
    QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
    QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
    QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
    getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
    getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
    getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
    getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
    accessQueueMisc_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueMisc_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueMisc_call_data : out  std_logic_vector(104 downto 0);
    accessQueueMisc_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueMisc_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueMisc_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueMisc_return_data : in   std_logic_vector(31 downto 0);
    accessQueueMisc_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(71 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
    setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(103 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(63 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(71 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
    getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
    getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
    getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
    getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(71 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 18)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 65)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal queue_type_buffer :  std_logic_vector(1 downto 0);
  signal queue_type_update_enable: Boolean;
  signal server_id_buffer :  std_logic_vector(7 downto 0);
  signal server_id_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(63 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_1669_start: Boolean;
  signal popFromQueue_CP_1669_symbol: Boolean;
  -- volatile/operator module components. 
  component getQueuePointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLockPointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessQueueMisc is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock_address_pointer : in  std_logic_vector(63 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_data : out  std_logic_vector(135 downto 0);
      accessMemoryLdStub_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryLdStub_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
      accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      buf_base_addr : in  std_logic_vector(63 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(63 downto 0);
      accessQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_call_data : out  std_logic_vector(168 downto 0);
      accessQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_return_data : in   std_logic_vector(63 downto 0);
      accessQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      queue_length : out  std_logic_vector(31 downto 0);
      accessQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueLength_call_data : out  std_logic_vector(104 downto 0);
      accessQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueLength_return_data : in   std_logic_vector(31 downto 0);
      accessQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueBufPointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
      accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock_address_pointer : in  std_logic_vector(63 downto 0);
      accessMemoryByte_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByte_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByte_call_data : out  std_logic_vector(144 downto 0);
      accessMemoryByte_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryByte_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByte_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByte_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByte_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1208_call_req_0 : boolean;
  signal call_stmt_1208_call_ack_0 : boolean;
  signal call_stmt_1208_call_req_1 : boolean;
  signal call_stmt_1208_call_ack_1 : boolean;
  signal call_stmt_1216_call_req_0 : boolean;
  signal call_stmt_1216_call_ack_0 : boolean;
  signal call_stmt_1216_call_req_1 : boolean;
  signal call_stmt_1216_call_ack_1 : boolean;
  signal call_stmt_1226_call_req_0 : boolean;
  signal call_stmt_1226_call_ack_0 : boolean;
  signal call_stmt_1226_call_req_1 : boolean;
  signal call_stmt_1226_call_ack_1 : boolean;
  signal call_stmt_1231_call_req_0 : boolean;
  signal call_stmt_1231_call_ack_0 : boolean;
  signal call_stmt_1231_call_req_1 : boolean;
  signal call_stmt_1231_call_ack_1 : boolean;
  signal call_stmt_1237_call_req_0 : boolean;
  signal call_stmt_1237_call_ack_0 : boolean;
  signal call_stmt_1237_call_req_1 : boolean;
  signal call_stmt_1237_call_ack_1 : boolean;
  signal call_stmt_1241_call_req_0 : boolean;
  signal call_stmt_1241_call_ack_0 : boolean;
  signal call_stmt_1241_call_req_1 : boolean;
  signal call_stmt_1241_call_ack_1 : boolean;
  signal call_stmt_1245_call_req_0 : boolean;
  signal call_stmt_1245_call_ack_0 : boolean;
  signal call_stmt_1245_call_req_1 : boolean;
  signal call_stmt_1245_call_ack_1 : boolean;
  signal CONCAT_u16_u32_1266_inst_req_0 : boolean;
  signal CONCAT_u16_u32_1266_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_1266_inst_req_1 : boolean;
  signal CONCAT_u16_u32_1266_inst_ack_1 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_req_0 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_ack_0 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_req_1 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_ack_1 : boolean;
  signal call_stmt_1288_call_req_0 : boolean;
  signal call_stmt_1288_call_ack_0 : boolean;
  signal call_stmt_1288_call_req_1 : boolean;
  signal call_stmt_1288_call_ack_1 : boolean;
  signal call_stmt_1294_call_req_0 : boolean;
  signal call_stmt_1294_call_ack_0 : boolean;
  signal call_stmt_1294_call_req_1 : boolean;
  signal call_stmt_1294_call_ack_1 : boolean;
  signal call_stmt_1300_call_req_0 : boolean;
  signal call_stmt_1300_call_ack_0 : boolean;
  signal call_stmt_1300_call_req_1 : boolean;
  signal call_stmt_1300_call_ack_1 : boolean;
  signal call_stmt_1308_call_req_0 : boolean;
  signal call_stmt_1308_call_ack_0 : boolean;
  signal call_stmt_1308_call_req_1 : boolean;
  signal call_stmt_1308_call_ack_1 : boolean;
  signal CONCAT_u16_u32_1325_inst_req_0 : boolean;
  signal CONCAT_u16_u32_1325_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_1325_inst_req_1 : boolean;
  signal CONCAT_u16_u32_1325_inst_ack_1 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_req_0 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_ack_0 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_req_1 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_ack_1 : boolean;
  signal call_stmt_1331_call_req_0 : boolean;
  signal call_stmt_1331_call_ack_0 : boolean;
  signal call_stmt_1331_call_req_1 : boolean;
  signal call_stmt_1331_call_ack_1 : boolean;
  signal W_status_1332_inst_req_0 : boolean;
  signal W_status_1332_inst_ack_0 : boolean;
  signal W_status_1332_inst_req_1 : boolean;
  signal W_status_1332_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 18) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(9 downto 8) <= queue_type;
  queue_type_buffer <= in_buffer_data_out(9 downto 8);
  in_buffer_data_in(17 downto 10) <= server_id;
  server_id_buffer <= in_buffer_data_out(17 downto 10);
  in_buffer_data_in(tag_length + 17 downto 18) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 17 downto 18);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_1669_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 65) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(64 downto 64) <= status_buffer;
  status <= out_buffer_data_out(64 downto 64);
  out_buffer_data_in(tag_length + 64 downto 65) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 64 downto 65);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_1669_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_1669_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_1669_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_1669: Block -- control-path 
    signal popFromQueue_CP_1669_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_1669_elements(0) <= popFromQueue_CP_1669_start;
    popFromQueue_CP_1669_symbol <= popFromQueue_CP_1669_elements(39);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1208/$entry
      -- CP-element group 0: 	 call_stmt_1208/call_stmt_1208_sample_start_
      -- CP-element group 0: 	 call_stmt_1208/call_stmt_1208_update_start_
      -- CP-element group 0: 	 call_stmt_1208/call_stmt_1208_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1208/call_stmt_1208_Sample/crr
      -- CP-element group 0: 	 call_stmt_1208/call_stmt_1208_Update/$entry
      -- CP-element group 0: 	 call_stmt_1208/call_stmt_1208_Update/ccr
      -- 
    ccr_1687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(0), ack => call_stmt_1208_call_req_1); -- 
    crr_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(0), ack => call_stmt_1208_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1208/call_stmt_1208_sample_completed_
      -- CP-element group 1: 	 call_stmt_1208/call_stmt_1208_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1208/call_stmt_1208_Sample/cra
      -- 
    cra_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1208_call_ack_0, ack => popFromQueue_CP_1669_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_1208/$exit
      -- CP-element group 2: 	 call_stmt_1208/call_stmt_1208_update_completed_
      -- CP-element group 2: 	 call_stmt_1208/call_stmt_1208_Update/$exit
      -- CP-element group 2: 	 call_stmt_1208/call_stmt_1208_Update/cca
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/$entry
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_sample_start_
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_update_start_
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Sample/crr
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Update/$entry
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Update/ccr
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_update_start_
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Update/$entry
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Update/ccr
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_update_start_
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Update/$entry
      -- CP-element group 2: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Update/ccr
      -- 
    cca_1688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1208_call_ack_1, ack => popFromQueue_CP_1669_elements(2)); -- 
    crr_1699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(2), ack => call_stmt_1216_call_req_0); -- 
    ccr_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(2), ack => call_stmt_1216_call_req_1); -- 
    ccr_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(2), ack => call_stmt_1226_call_req_1); -- 
    ccr_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(2), ack => call_stmt_1231_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_sample_completed_
      -- CP-element group 3: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Sample/cra
      -- 
    cra_1700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1216_call_ack_0, ack => popFromQueue_CP_1669_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_update_completed_
      -- CP-element group 4: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Update/$exit
      -- CP-element group 4: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1216_Update/cca
      -- CP-element group 4: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_sample_start_
      -- CP-element group 4: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Sample/crr
      -- 
    cca_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1216_call_ack_1, ack => popFromQueue_CP_1669_elements(4)); -- 
    crr_1713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(4), ack => call_stmt_1226_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_sample_completed_
      -- CP-element group 5: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Sample/$exit
      -- CP-element group 5: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Sample/cra
      -- 
    cra_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1226_call_ack_0, ack => popFromQueue_CP_1669_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_update_completed_
      -- CP-element group 6: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Update/$exit
      -- CP-element group 6: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1226_Update/cca
      -- 
    cca_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1226_call_ack_1, ack => popFromQueue_CP_1669_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_sample_start_
      -- CP-element group 7: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Sample/$entry
      -- CP-element group 7: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Sample/crr
      -- 
    crr_1727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(7), ack => call_stmt_1231_call_req_0); -- 
    popFromQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "popFromQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1669_elements(4) & popFromQueue_CP_1669_elements(6);
      gj_popFromQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1669_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_sample_completed_
      -- CP-element group 8: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Sample/$exit
      -- CP-element group 8: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Sample/cra
      -- 
    cra_1728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1231_call_ack_0, ack => popFromQueue_CP_1669_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	18 
    -- CP-element group 9:  members (20) 
      -- CP-element group 9: 	 call_stmt_1216_to_call_stmt_1231/$exit
      -- CP-element group 9: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_update_completed_
      -- CP-element group 9: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Update/$exit
      -- CP-element group 9: 	 call_stmt_1216_to_call_stmt_1231/call_stmt_1231_Update/cca
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/$entry
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_sample_start_
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_update_start_
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Sample/$entry
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Sample/crr
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Update/$entry
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Update/ccr
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_update_start_
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Update/$entry
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Update/ccr
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_update_start_
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Update/$entry
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Update/ccr
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_update_start_
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Update/$entry
      -- CP-element group 9: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Update/cr
      -- 
    cca_1733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1231_call_ack_1, ack => popFromQueue_CP_1669_elements(9)); -- 
    crr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(9), ack => call_stmt_1237_call_req_0); -- 
    ccr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(9), ack => call_stmt_1237_call_req_1); -- 
    ccr_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(9), ack => call_stmt_1241_call_req_1); -- 
    ccr_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(9), ack => call_stmt_1245_call_req_1); -- 
    cr_1791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(9), ack => CONCAT_u16_u32_1266_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_sample_completed_
      -- CP-element group 10: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Sample/$exit
      -- CP-element group 10: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Sample/cra
      -- 
    cra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1237_call_ack_0, ack => popFromQueue_CP_1669_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	16 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_update_completed_
      -- CP-element group 11: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Update/$exit
      -- CP-element group 11: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1237_Update/cca
      -- CP-element group 11: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_sample_start_
      -- CP-element group 11: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Sample/$entry
      -- CP-element group 11: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Sample/crr
      -- 
    cca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1237_call_ack_1, ack => popFromQueue_CP_1669_elements(11)); -- 
    crr_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(11), ack => call_stmt_1241_call_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_sample_completed_
      -- CP-element group 12: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Sample/$exit
      -- CP-element group 12: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Sample/cra
      -- 
    cra_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1241_call_ack_0, ack => popFromQueue_CP_1669_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_update_completed_
      -- CP-element group 13: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Update/$exit
      -- CP-element group 13: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1241_Update/cca
      -- CP-element group 13: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_sample_start_
      -- CP-element group 13: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Sample/$entry
      -- CP-element group 13: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Sample/crr
      -- 
    cca_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1241_call_ack_1, ack => popFromQueue_CP_1669_elements(13)); -- 
    crr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(13), ack => call_stmt_1245_call_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_sample_completed_
      -- CP-element group 14: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Sample/$exit
      -- CP-element group 14: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Sample/cra
      -- 
    cra_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1245_call_ack_0, ack => popFromQueue_CP_1669_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	19 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_update_completed_
      -- CP-element group 15: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Update/$exit
      -- CP-element group 15: 	 call_stmt_1237_to_assign_stmt_1267/call_stmt_1245_Update/cca
      -- 
    cca_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1245_call_ack_1, ack => popFromQueue_CP_1669_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_sample_start_
      -- CP-element group 16: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Sample/$entry
      -- CP-element group 16: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Sample/rr
      -- 
    rr_1786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(16), ack => CONCAT_u16_u32_1266_inst_req_0); -- 
    popFromQueue_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1669_elements(11) & popFromQueue_CP_1669_elements(15);
      gj_popFromQueue_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1669_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_sample_completed_
      -- CP-element group 17: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Sample/$exit
      -- CP-element group 17: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Sample/ra
      -- 
    ra_1787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1266_inst_ack_0, ack => popFromQueue_CP_1669_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	9 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_update_completed_
      -- CP-element group 18: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Update/$exit
      -- CP-element group 18: 	 call_stmt_1237_to_assign_stmt_1267/CONCAT_u16_u32_1266_Update/ca
      -- 
    ca_1792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1266_inst_ack_1, ack => popFromQueue_CP_1669_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_sample_start_
      -- CP-element group 19: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Sample/req
      -- 
    req_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(19), ack => WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_req_0); -- 
    popFromQueue_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1669_elements(15) & popFromQueue_CP_1669_elements(18);
      gj_popFromQueue_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1669_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_sample_completed_
      -- CP-element group 20: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_update_start_
      -- CP-element group 20: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Sample/ack
      -- CP-element group 20: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Update/$entry
      -- CP-element group 20: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Update/req
      -- 
    ack_1801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_ack_0, ack => popFromQueue_CP_1669_elements(20)); -- 
    req_1805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(20), ack => WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	27 
    -- CP-element group 21: 	29 
    -- CP-element group 21: 	30 
    -- CP-element group 21: 	31 
    -- CP-element group 21:  members (26) 
      -- CP-element group 21: 	 call_stmt_1237_to_assign_stmt_1267/$exit
      -- CP-element group 21: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_update_completed_
      -- CP-element group 21: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Update/$exit
      -- CP-element group 21: 	 call_stmt_1237_to_assign_stmt_1267/WPIPE_QUEUE_MONITOR_SIGNAL_1252_Update/ack
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_sample_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_update_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Sample/crr
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Update/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Update/ccr
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_update_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Update/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Update/ccr
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_update_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Update/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Update/ccr
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_update_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Update/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Update/ccr
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_sample_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_update_start_
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Sample/rr
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Update/$entry
      -- CP-element group 21: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Update/cr
      -- 
    ack_1806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_ack_1, ack => popFromQueue_CP_1669_elements(21)); -- 
    crr_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => call_stmt_1288_call_req_0); -- 
    ccr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => call_stmt_1288_call_req_1); -- 
    ccr_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => call_stmt_1294_call_req_1); -- 
    ccr_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => call_stmt_1300_call_req_1); -- 
    ccr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => call_stmt_1308_call_req_1); -- 
    rr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => CONCAT_u16_u32_1325_inst_req_0); -- 
    cr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(21), ack => CONCAT_u16_u32_1325_inst_req_1); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_sample_completed_
      -- CP-element group 22: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Sample/$exit
      -- CP-element group 22: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Sample/cra
      -- 
    cra_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1288_call_ack_0, ack => popFromQueue_CP_1669_elements(22)); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_update_completed_
      -- CP-element group 23: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Update/$exit
      -- CP-element group 23: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1288_Update/cca
      -- CP-element group 23: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_sample_start_
      -- CP-element group 23: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Sample/crr
      -- 
    cca_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1288_call_ack_1, ack => popFromQueue_CP_1669_elements(23)); -- 
    crr_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(23), ack => call_stmt_1294_call_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_sample_completed_
      -- CP-element group 24: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Sample/cra
      -- 
    cra_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1294_call_ack_0, ack => popFromQueue_CP_1669_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	21 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_update_completed_
      -- CP-element group 25: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Update/$exit
      -- CP-element group 25: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1294_Update/cca
      -- CP-element group 25: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_sample_start_
      -- CP-element group 25: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Sample/crr
      -- 
    cca_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1294_call_ack_1, ack => popFromQueue_CP_1669_elements(25)); -- 
    crr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(25), ack => call_stmt_1300_call_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_sample_completed_
      -- CP-element group 26: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Sample/$exit
      -- CP-element group 26: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Sample/cra
      -- 
    cra_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1300_call_ack_0, ack => popFromQueue_CP_1669_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	21 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_update_completed_
      -- CP-element group 27: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Update/$exit
      -- CP-element group 27: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1300_Update/cca
      -- CP-element group 27: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_sample_start_
      -- CP-element group 27: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Sample/crr
      -- 
    cca_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1300_call_ack_1, ack => popFromQueue_CP_1669_elements(27)); -- 
    crr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(27), ack => call_stmt_1308_call_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_sample_completed_
      -- CP-element group 28: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Sample/cra
      -- 
    cra_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1308_call_ack_0, ack => popFromQueue_CP_1669_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	21 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_update_completed_
      -- CP-element group 29: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Update/$exit
      -- CP-element group 29: 	 assign_stmt_1275_to_assign_stmt_1326/call_stmt_1308_Update/cca
      -- 
    cca_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1308_call_ack_1, ack => popFromQueue_CP_1669_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	21 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_sample_completed_
      -- CP-element group 30: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Sample/$exit
      -- CP-element group 30: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Sample/ra
      -- 
    ra_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1325_inst_ack_0, ack => popFromQueue_CP_1669_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	21 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_update_completed_
      -- CP-element group 31: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Update/$exit
      -- CP-element group 31: 	 assign_stmt_1275_to_assign_stmt_1326/CONCAT_u16_u32_1325_Update/ca
      -- CP-element group 31: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_sample_start_
      -- CP-element group 31: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Sample/$entry
      -- CP-element group 31: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Sample/req
      -- 
    ca_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1325_inst_ack_1, ack => popFromQueue_CP_1669_elements(31)); -- 
    req_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(31), ack => WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_sample_completed_
      -- CP-element group 32: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_update_start_
      -- CP-element group 32: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Sample/ack
      -- CP-element group 32: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Update/$entry
      -- CP-element group 32: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Update/req
      -- 
    ack_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_ack_0, ack => popFromQueue_CP_1669_elements(32)); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(32), ack => WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_update_completed_
      -- CP-element group 33: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Update/$exit
      -- CP-element group 33: 	 assign_stmt_1275_to_assign_stmt_1326/WPIPE_QUEUE_MONITOR_SIGNAL_1310_Update/ack
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_ack_1, ack => popFromQueue_CP_1669_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34:  members (14) 
      -- CP-element group 34: 	 assign_stmt_1275_to_assign_stmt_1326/$exit
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/$entry
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_sample_start_
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_update_start_
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Sample/$entry
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Sample/crr
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Update/$entry
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Update/ccr
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_sample_start_
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_update_start_
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Sample/$entry
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Sample/req
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Update/$entry
      -- CP-element group 34: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Update/req
      -- 
    crr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(34), ack => call_stmt_1331_call_req_0); -- 
    ccr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(34), ack => call_stmt_1331_call_req_1); -- 
    req_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(34), ack => W_status_1332_inst_req_0); -- 
    req_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1669_elements(34), ack => W_status_1332_inst_req_1); -- 
    popFromQueue_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1669_elements(29) & popFromQueue_CP_1669_elements(33);
      gj_popFromQueue_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1669_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_sample_completed_
      -- CP-element group 35: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Sample/$exit
      -- CP-element group 35: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Sample/cra
      -- 
    cra_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1331_call_ack_0, ack => popFromQueue_CP_1669_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	39 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_update_completed_
      -- CP-element group 36: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Update/$exit
      -- CP-element group 36: 	 call_stmt_1331_to_assign_stmt_1334/call_stmt_1331_Update/cca
      -- 
    cca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1331_call_ack_1, ack => popFromQueue_CP_1669_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_sample_completed_
      -- CP-element group 37: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Sample/$exit
      -- CP-element group 37: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Sample/ack
      -- 
    ack_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1332_inst_ack_0, ack => popFromQueue_CP_1669_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_update_completed_
      -- CP-element group 38: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Update/$exit
      -- CP-element group 38: 	 call_stmt_1331_to_assign_stmt_1334/assign_stmt_1334_Update/ack
      -- 
    ack_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1332_inst_ack_1, ack => popFromQueue_CP_1669_elements(38)); -- 
    -- CP-element group 39:  join  transition  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	36 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 $exit
      -- CP-element group 39: 	 call_stmt_1331_to_assign_stmt_1334/$exit
      -- 
    popFromQueue_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1669_elements(36) & popFromQueue_CP_1669_elements(38);
      gj_popFromQueue_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1669_elements(39), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1281_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1266_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1325_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u4_u8_1256_wire : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_1314_wire : std_logic_vector(7 downto 0);
    signal CONCAT_u8_u16_1259_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_1264_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_1319_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_1324_wire : std_logic_vector(15 downto 0);
    signal R_POPQ_1313_wire_constant : std_logic_vector(3 downto 0);
    signal R_PREPOPQ_1255_wire_constant : std_logic_vector(3 downto 0);
    signal R_READMEM_1211_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u32_u32_1273_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1307_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1317_wire : std_logic_vector(31 downto 0);
    signal konst_1219_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1248_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1272_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1278_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1280_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1316_wire_constant : std_logic_vector(31 downto 0);
    signal lock_n_1221 : std_logic_vector(0 downto 0);
    signal m_ok_1231 : std_logic_vector(0 downto 0);
    signal misc_1216 : std_logic_vector(31 downto 0);
    signal next_ri_1283 : std_logic_vector(31 downto 0);
    signal q_base_address_1208 : std_logic_vector(63 downto 0);
    signal q_buf_address_1288 : std_logic_vector(63 downto 0);
    signal q_empty_1250 : std_logic_vector(0 downto 0);
    signal q_lock_address_1226 : std_logic_vector(63 downto 0);
    signal queue_length_1241 : std_logic_vector(31 downto 0);
    signal read_index_1237 : std_logic_vector(31 downto 0);
    signal round_off_1275 : std_logic_vector(0 downto 0);
    signal total_msgs_1245 : std_logic_vector(31 downto 0);
    signal type_cast_1214_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1254_wire : std_logic_vector(3 downto 0);
    signal type_cast_1258_wire : std_logic_vector(7 downto 0);
    signal type_cast_1261_wire : std_logic_vector(7 downto 0);
    signal type_cast_1263_wire : std_logic_vector(7 downto 0);
    signal type_cast_1306_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1312_wire : std_logic_vector(3 downto 0);
    signal type_cast_1318_wire : std_logic_vector(7 downto 0);
    signal type_cast_1321_wire : std_logic_vector(7 downto 0);
    signal type_cast_1323_wire : std_logic_vector(7 downto 0);
    signal write_index_1237 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_POPQ_1313_wire_constant <= "0001";
    R_PREPOPQ_1255_wire_constant <= "0011";
    R_READMEM_1211_wire_constant <= "1";
    konst_1219_wire_constant <= "00000000000000000000000000000000";
    konst_1248_wire_constant <= "00000000000000000000000000000000";
    konst_1272_wire_constant <= "00000000000000000000000000000001";
    konst_1278_wire_constant <= "00000000000000000000000000000000";
    konst_1280_wire_constant <= "00000000000000000000000000000001";
    konst_1316_wire_constant <= "00000000000000000000000000000001";
    type_cast_1214_wire_constant <= "00000000000000000000000000000000";
    type_cast_1306_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_1282_inst
    next_ri_1283 <= konst_1278_wire_constant when (round_off_1275(0) /=  '0') else ADD_u32_u32_1281_wire;
    W_status_1332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_1332_inst_req_0;
      W_status_1332_inst_ack_0<= wack(0);
      rreq(0) <= W_status_1332_inst_req_1;
      W_status_1332_inst_ack_1<= rack(0);
      W_status_1332_inst : InterlockBuffer generic map ( -- 
        name => "W_status_1332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_empty_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1254_inst
    process(queue_type_buffer) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := queue_type_buffer(1 downto 0);
      type_cast_1254_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1258_inst
    process(total_msgs_1245) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := total_msgs_1245(7 downto 0);
      type_cast_1258_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1261_inst
    process(write_index_1237) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := write_index_1237(7 downto 0);
      type_cast_1261_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1263_inst
    process(read_index_1237) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := read_index_1237(7 downto 0);
      type_cast_1263_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1312_inst
    process(queue_type_buffer) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := queue_type_buffer(1 downto 0);
      type_cast_1312_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1318_inst
    process(SUB_u32_u32_1317_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u32_u32_1317_wire(7 downto 0);
      type_cast_1318_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1321_inst
    process(write_index_1237) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := write_index_1237(7 downto 0);
      type_cast_1321_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1323_inst
    process(next_ri_1283) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := next_ri_1283(7 downto 0);
      type_cast_1323_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator ADD_u32_u32_1281_inst
    ADD_u32_u32_1281_wire <= std_logic_vector(unsigned(read_index_1237) + unsigned(konst_1280_wire_constant));
    -- flow through binary operator BITSEL_u32_u1_1220_inst
    process(misc_1216) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(misc_1216, konst_1219_wire_constant, tmp_var);
      lock_n_1221 <= tmp_var; --
    end process;
    -- shared split operator group (2) : CONCAT_u16_u32_1266_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_1259_wire & CONCAT_u8_u16_1264_wire;
      CONCAT_u16_u32_1266_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  not q_empty_1250(0);
      reqL_unguarded(0) <= CONCAT_u16_u32_1266_inst_req_0;
      CONCAT_u16_u32_1266_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_1266_inst_req_1;
      CONCAT_u16_u32_1266_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : CONCAT_u16_u32_1325_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_1319_wire & CONCAT_u8_u16_1324_wire;
      CONCAT_u16_u32_1325_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  not q_empty_1250(0);
      reqL_unguarded(0) <= CONCAT_u16_u32_1325_inst_req_0;
      CONCAT_u16_u32_1325_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_1325_inst_req_1;
      CONCAT_u16_u32_1325_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- flow through binary operator CONCAT_u4_u8_1256_inst
    process(type_cast_1254_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1254_wire, R_PREPOPQ_1255_wire_constant, tmp_var);
      CONCAT_u4_u8_1256_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u8_1314_inst
    process(type_cast_1312_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1312_wire, R_POPQ_1313_wire_constant, tmp_var);
      CONCAT_u4_u8_1314_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_1259_inst
    process(CONCAT_u4_u8_1256_wire, type_cast_1258_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u8_1256_wire, type_cast_1258_wire, tmp_var);
      CONCAT_u8_u16_1259_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_1264_inst
    process(type_cast_1261_wire, type_cast_1263_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1261_wire, type_cast_1263_wire, tmp_var);
      CONCAT_u8_u16_1264_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_1319_inst
    process(CONCAT_u4_u8_1314_wire, type_cast_1318_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u8_1314_wire, type_cast_1318_wire, tmp_var);
      CONCAT_u8_u16_1319_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_1324_inst
    process(type_cast_1321_wire, type_cast_1323_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1321_wire, type_cast_1323_wire, tmp_var);
      CONCAT_u8_u16_1324_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_1249_inst
    process(total_msgs_1245) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(total_msgs_1245, konst_1248_wire_constant, tmp_var);
      q_empty_1250 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_1274_inst
    process(read_index_1237, SUB_u32_u32_1273_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(read_index_1237, SUB_u32_u32_1273_wire, tmp_var);
      round_off_1275 <= tmp_var; --
    end process;
    -- flow through binary operator SUB_u32_u32_1273_inst
    SUB_u32_u32_1273_wire <= std_logic_vector(unsigned(queue_length_1241) - unsigned(konst_1272_wire_constant));
    -- flow through binary operator SUB_u32_u32_1307_inst
    SUB_u32_u32_1307_wire <= std_logic_vector(unsigned(total_msgs_1245) - unsigned(type_cast_1306_wire_constant));
    -- flow through binary operator SUB_u32_u32_1317_inst
    SUB_u32_u32_1317_wire <= std_logic_vector(unsigned(total_msgs_1245) - unsigned(konst_1316_wire_constant));
    -- shared outport operator group (0) : WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_req_0;
      WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_req_1;
      update_req_unguarded(0) <= WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_req_1;
      WPIPE_QUEUE_MONITOR_SIGNAL_1310_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_QUEUE_MONITOR_SIGNAL_1252_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not q_empty_1250(0);
      guard_vector(1)  <=  not q_empty_1250(0);
      data_in <= CONCAT_u16_u32_1325_wire & CONCAT_u16_u32_1266_wire;
      QUEUE_MONITOR_SIGNAL_write_0_gI: SplitGuardInterface generic map(name => "QUEUE_MONITOR_SIGNAL_write_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      QUEUE_MONITOR_SIGNAL_write_0: OutputPortRevised -- 
        generic map ( name => "QUEUE_MONITOR_SIGNAL", data_width => 32, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => QUEUE_MONITOR_SIGNAL_pipe_write_req(0),
          oack => QUEUE_MONITOR_SIGNAL_pipe_write_ack(0),
          odata => QUEUE_MONITOR_SIGNAL_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1208_call 
    getQueuePointer_call_group_0: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1208_call_req_0;
      call_stmt_1208_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1208_call_req_1;
      call_stmt_1208_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointer_call_group_0_gI: SplitGuardInterface generic map(name => "getQueuePointer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= queue_type_buffer & server_id_buffer;
      q_base_address_1208 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 10,
        owidth => 10,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointer_call_reqs(0),
          ackR => getQueuePointer_call_acks(0),
          dataR => getQueuePointer_call_data(9 downto 0),
          tagR => getQueuePointer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointer_return_acks(0), -- cross-over
          ackL => getQueuePointer_return_reqs(0), -- cross-over
          dataL => getQueuePointer_return_data(63 downto 0),
          tagL => getQueuePointer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1216_call 
    accessQueueMisc_call_group_1: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1216_call_req_0;
      call_stmt_1216_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1216_call_req_1;
      call_stmt_1216_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueMisc_call_group_1_gI: SplitGuardInterface generic map(name => "accessQueueMisc_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_1211_wire_constant & q_base_address_1208 & type_cast_1214_wire_constant;
      misc_1216 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueMisc_call_reqs(0),
          ackR => accessQueueMisc_call_acks(0),
          dataR => accessQueueMisc_call_data(104 downto 0),
          tagR => accessQueueMisc_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueMisc_return_acks(0), -- cross-over
          ackL => accessQueueMisc_return_reqs(0), -- cross-over
          dataL => accessQueueMisc_return_data(31 downto 0),
          tagL => accessQueueMisc_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1226_call 
    getQueueLockPointer_call_group_2: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1226_call_req_0;
      call_stmt_1226_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1226_call_req_1;
      call_stmt_1226_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not lock_n_1221(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLockPointer_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueLockPointer_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= queue_type_buffer & server_id_buffer;
      q_lock_address_1226 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 10,
        owidth => 10,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLockPointer_call_reqs(0),
          ackR => getQueueLockPointer_call_acks(0),
          dataR => getQueueLockPointer_call_data(9 downto 0),
          tagR => getQueueLockPointer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLockPointer_return_acks(0), -- cross-over
          ackL => getQueueLockPointer_return_reqs(0), -- cross-over
          dataL => getQueueLockPointer_return_data(63 downto 0),
          tagL => getQueueLockPointer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1231_call 
    acquireLock_call_group_3: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1231_call_req_0;
      call_stmt_1231_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1231_call_req_1;
      call_stmt_1231_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not lock_n_1221(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_3_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_lock_address_1226;
      m_ok_1231 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(71 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1237_call 
    getQueuePointers_call_group_4: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1237_call_req_0;
      call_stmt_1237_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1237_call_req_1;
      call_stmt_1237_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_4_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1208;
      write_index_1237 <= data_out(63 downto 32);
      read_index_1237 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(71 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1241_call 
    getQueueLength_call_group_5: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1241_call_req_0;
      call_stmt_1241_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1241_call_req_1;
      call_stmt_1241_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_5_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1208;
      queue_length_1241 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(71 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1245_call 
    getTotalMessages_call_group_6: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1245_call_req_0;
      call_stmt_1245_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1245_call_req_1;
      call_stmt_1245_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_6_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1208;
      total_msgs_1245 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(71 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1288_call 
    getQueueBufPointer_call_group_7: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1288_call_req_0;
      call_stmt_1288_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1288_call_req_1;
      call_stmt_1288_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1250(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueBufPointer_call_group_7_gI: SplitGuardInterface generic map(name => "getQueueBufPointer_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= queue_type_buffer & server_id_buffer;
      q_buf_address_1288 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 10,
        owidth => 10,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueBufPointer_call_reqs(0),
          ackR => getQueueBufPointer_call_acks(0),
          dataR => getQueueBufPointer_call_data(9 downto 0),
          tagR => getQueueBufPointer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueBufPointer_return_acks(0), -- cross-over
          ackL => getQueueBufPointer_return_reqs(0), -- cross-over
          dataL => getQueueBufPointer_return_data(63 downto 0),
          tagL => getQueueBufPointer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_1294_call 
    getQueueElement_call_group_8: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1294_call_req_0;
      call_stmt_1294_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1294_call_req_1;
      call_stmt_1294_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1250(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_8_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_buf_address_1288 & read_index_1237;
      q_r_data_buffer <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(103 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(63 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- shared call operator group (9) : call_stmt_1300_call 
    setQueuePointers_call_group_9: Block -- 
      signal data_in: std_logic_vector(135 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1300_call_req_0;
      call_stmt_1300_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1300_call_req_1;
      call_stmt_1300_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1250(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_9_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1208 & write_index_1237 & next_ri_1283;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 136,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(135 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 9
    -- shared call operator group (10) : call_stmt_1308_call 
    setTotalMessages_call_group_10: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1308_call_req_0;
      call_stmt_1308_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1308_call_req_1;
      call_stmt_1308_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1250(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setTotalMessages_call_group_10_gI: SplitGuardInterface generic map(name => "setTotalMessages_call_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1208 & SUB_u32_u32_1307_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setTotalMessages_call_reqs(0),
          ackR => setTotalMessages_call_acks(0),
          dataR => setTotalMessages_call_data(103 downto 0),
          tagR => setTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setTotalMessages_return_acks(0), -- cross-over
          ackL => setTotalMessages_return_reqs(0), -- cross-over
          tagL => setTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 10
    -- shared call operator group (11) : call_stmt_1331_call 
    releaseLock_call_group_11: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1331_call_req_0;
      call_stmt_1331_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1331_call_req_1;
      call_stmt_1331_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not lock_n_1221(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_11_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_lock_address_1226;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(71 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 11
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    rx_buffer_pointer : in  std_logic_vector(63 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(7 downto 0);
    S_NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(7 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    incrementNumberOfPacketsReceived_call_reqs : out  std_logic_vector(0 downto 0);
    incrementNumberOfPacketsReceived_call_acks : in   std_logic_vector(0 downto 0);
    incrementNumberOfPacketsReceived_call_tag  :  out  std_logic_vector(0 downto 0);
    incrementNumberOfPacketsReceived_return_reqs : out  std_logic_vector(0 downto 0);
    incrementNumberOfPacketsReceived_return_acks : in   std_logic_vector(0 downto 0);
    incrementNumberOfPacketsReceived_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal rx_buffer_pointer_buffer :  std_logic_vector(63 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_2805_start: Boolean;
  signal populateRxQueue_CP_2805_symbol: Boolean;
  -- volatile/operator module components. 
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_w_data : in  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(167 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(9 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  component incrementNumberOfPacketsReceived is -- 
    generic (tag_length : integer); 
    port ( -- 
      incrementRegister_call_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_call_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_call_data : out  std_logic_vector(7 downto 0);
      incrementRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementRegister_return_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_return_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_return_data : in   std_logic_vector(31 downto 0);
      incrementRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1773_call_ack_1 : boolean;
  signal call_stmt_1775_call_ack_1 : boolean;
  signal call_stmt_1794_call_req_0 : boolean;
  signal call_stmt_1773_call_req_1 : boolean;
  signal call_stmt_1773_call_ack_0 : boolean;
  signal call_stmt_1773_call_req_0 : boolean;
  signal call_stmt_1775_call_req_1 : boolean;
  signal call_stmt_1794_call_ack_1 : boolean;
  signal call_stmt_1775_call_req_0 : boolean;
  signal call_stmt_1794_call_ack_0 : boolean;
  signal call_stmt_1775_call_ack_0 : boolean;
  signal if_stmt_1789_branch_ack_1 : boolean;
  signal call_stmt_1794_call_req_1 : boolean;
  signal AND_u8_u8_1784_inst_ack_1 : boolean;
  signal AND_u8_u8_1784_inst_req_1 : boolean;
  signal AND_u8_u8_1784_inst_ack_0 : boolean;
  signal if_stmt_1789_branch_ack_0 : boolean;
  signal if_stmt_1789_branch_req_0 : boolean;
  signal AND_u8_u8_1784_inst_req_0 : boolean;
  signal if_stmt_1795_branch_req_0 : boolean;
  signal if_stmt_1795_branch_ack_1 : boolean;
  signal if_stmt_1795_branch_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_ack_1 : boolean;
  signal AND_u8_u8_1763_inst_req_0 : boolean;
  signal AND_u8_u8_1763_inst_ack_0 : boolean;
  signal AND_u8_u8_1763_inst_req_1 : boolean;
  signal AND_u8_u8_1763_inst_ack_1 : boolean;
  signal phi_stmt_1754_req_0 : boolean;
  signal n_q_index_1785_1764_buf_req_0 : boolean;
  signal n_q_index_1785_1764_buf_ack_0 : boolean;
  signal n_q_index_1785_1764_buf_req_1 : boolean;
  signal n_q_index_1785_1764_buf_ack_1 : boolean;
  signal phi_stmt_1754_req_1 : boolean;
  signal phi_stmt_1754_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_2805_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_2805_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_2805_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_2805_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_2805: Block -- control-path 
    signal populateRxQueue_CP_2805_elements: BooleanArray(26 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_2805_elements(0) <= populateRxQueue_CP_2805_start;
    populateRxQueue_CP_2805_symbol <= populateRxQueue_CP_2805_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	18 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 branch_block_stmt_1752/branch_block_stmt_1752__entry__
      -- CP-element group 0: 	 branch_block_stmt_1752/merge_stmt_1753__entry__
      -- CP-element group 0: 	 branch_block_stmt_1752/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1752/merge_stmt_1753_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	15 
    -- CP-element group 1: 	17 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1752/if_stmt_1789__exit__
      -- CP-element group 1: 	 branch_block_stmt_1752/branch_block_stmt_1752__exit__
      -- CP-element group 1: 	 branch_block_stmt_1752/$exit
      -- CP-element group 1: 	 $exit
      -- 
    populateRxQueue_CP_2805_elements(1) <= OrReduce(populateRxQueue_CP_2805_elements(15) & populateRxQueue_CP_2805_elements(17));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	26 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Sample/cra
      -- CP-element group 2: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_sample_completed_
      -- 
    cra_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1773_call_ack_0, ack => populateRxQueue_CP_2805_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	26 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	8 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_update_completed_
      -- 
    cca_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1773_call_ack_1, ack => populateRxQueue_CP_2805_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Sample/cra
      -- CP-element group 4: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Sample/$exit
      -- 
    cra_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1775_call_ack_0, ack => populateRxQueue_CP_2805_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	26 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	9 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Update/cca
      -- CP-element group 5: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_update_completed_
      -- 
    cca_2849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1775_call_ack_1, ack => populateRxQueue_CP_2805_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	26 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Sample/ra
      -- 
    ra_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u8_u8_1784_inst_ack_0, ack => populateRxQueue_CP_2805_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	26 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Update/$exit
      -- 
    ca_2863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u8_u8_1784_inst_ack_1, ack => populateRxQueue_CP_2805_elements(7)); -- 
    -- CP-element group 8:  transition  output  delay-element  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	4 
    -- CP-element group 8:  members (4) 
      -- CP-element group 8: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Sample/crr
      -- CP-element group 8: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_call_stmt_1775_delay
      -- CP-element group 8: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Sample/$entry
      -- 
    crr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(8), ack => call_stmt_1775_call_req_0); -- 
    -- Element group populateRxQueue_CP_2805_elements(8) is a control-delay.
    cp_element_8_delay: control_delay_element  generic map(name => " 8_delay", delay_value => 1)  port map(req => populateRxQueue_CP_2805_elements(3), ack => populateRxQueue_CP_2805_elements(8), clk => clk, reset =>reset);
    -- CP-element group 9:  branch  join  transition  place  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	5 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (22) 
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/NOT_u1_u1_1791_place
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_else_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/$exit
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789__entry__
      -- CP-element group 9: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785__exit__
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/$exit
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/SplitProtocol/$entry
      -- CP-element group 9: 	 branch_block_stmt_1752/if_stmt_1789_eval_test/NOT_u1_u1_1791/$exit
      -- 
    branch_req_2888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(9), ack => if_stmt_1789_branch_req_0); -- 
    populateRxQueue_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "populateRxQueue_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_2805_elements(5) & populateRxQueue_CP_2805_elements(7);
      gj_populateRxQueue_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_2805_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 branch_block_stmt_1752/if_stmt_1789_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Sample/crr
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1752/if_stmt_1789_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Update/ccr
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794/$entry
      -- CP-element group 10: 	 branch_block_stmt_1752/call_stmt_1794__entry__
      -- 
    if_choice_transition_2893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1789_branch_ack_1, ack => populateRxQueue_CP_2805_elements(10)); -- 
    crr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(10), ack => call_stmt_1794_call_req_0); -- 
    ccr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(10), ack => call_stmt_1794_call_req_1); -- 
    -- CP-element group 11:  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	16 
    -- CP-element group 11:  members (7) 
      -- CP-element group 11: 	 branch_block_stmt_1752/if_stmt_1789_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_1752/if_stmt_1789_else_link/else_choice_transition
      -- CP-element group 11: 	 branch_block_stmt_1752/assign_stmt_1804__entry__
      -- CP-element group 11: 	 branch_block_stmt_1752/assign_stmt_1804/$entry
      -- CP-element group 11: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Sample/req
      -- 
    else_choice_transition_2897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1789_branch_ack_0, ack => populateRxQueue_CP_2805_elements(11)); -- 
    req_2968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(11), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Sample/cra
      -- CP-element group 12: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_sample_completed_
      -- 
    cra_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1794_call_ack_0, ack => populateRxQueue_CP_2805_elements(12)); -- 
    -- CP-element group 13:  branch  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (27) 
      -- CP-element group 13: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Update/cca
      -- CP-element group 13: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/call_stmt_1794/call_stmt_1794_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_dead_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/call_stmt_1794/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/EQ_u1_u1_1798_inputs/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/EQ_u1_u1_1798_inputs/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795__entry__
      -- CP-element group 13: 	 branch_block_stmt_1752/call_stmt_1794__exit__
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/EQ_u1_u1_1798/SplitProtocol/Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_eval_test/branch_req
      -- CP-element group 13: 	 branch_block_stmt_1752/EQ_u1_u1_1798_place
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_if_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_1752/if_stmt_1795_else_link/$entry
      -- 
    cca_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1794_call_ack_1, ack => populateRxQueue_CP_2805_elements(13)); -- 
    branch_req_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(13), ack => if_stmt_1795_branch_req_0); -- 
    -- CP-element group 14:  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	22 
    -- CP-element group 14: 	23 
    -- CP-element group 14:  members (11) 
      -- CP-element group 14: 	 branch_block_stmt_1752/if_stmt_1795_if_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_1752/if_stmt_1795_if_link/if_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/$entry
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/$entry
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Sample/req
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Update/req
      -- 
    if_choice_transition_2950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1795_branch_ack_1, ack => populateRxQueue_CP_2805_elements(14)); -- 
    req_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(14), ack => n_q_index_1785_1764_buf_req_0); -- 
    req_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(14), ack => n_q_index_1785_1764_buf_req_1); -- 
    -- CP-element group 15:  merge  transition  place  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	1 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1752/if_stmt_1795__exit__
      -- CP-element group 15: 	 branch_block_stmt_1752/if_stmt_1795_else_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_1752/if_stmt_1795_else_link/else_choice_transition
      -- 
    else_choice_transition_2954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1795_branch_ack_0, ack => populateRxQueue_CP_2805_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Sample/ack
      -- CP-element group 16: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Update/req
      -- 
    ack_2969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_ack_0, ack => populateRxQueue_CP_2805_elements(16)); -- 
    req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(16), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_req_1); -- 
    -- CP-element group 17:  transition  place  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	1 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1752/assign_stmt_1804__exit__
      -- CP-element group 17: 	 branch_block_stmt_1752/assign_stmt_1804/$exit
      -- CP-element group 17: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1752/assign_stmt_1804/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_Update/ack
      -- 
    ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_ack_1, ack => populateRxQueue_CP_2805_elements(17)); -- 
    -- CP-element group 18:  join  fork  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (71) 
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Sample/req
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Update/req
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/ADD_u8_u8_1758_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756/Update/ack
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/ADD_u8_u8_1758/SplitProtocol/Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Sample/req
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Update/req
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SUB_u32_u32_1761_inputs/RPIPE_S_NUMBER_OF_SERVERS_1759/Update/ack
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SUB_u32_u32_1761/SplitProtocol/Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/AND_u8_u8_1763_inputs/type_cast_1762/SplitProtocol/Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Update/cr
      -- 
    cr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(18), ack => AND_u8_u8_1763_inst_req_1); -- 
    rr_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(18), ack => AND_u8_u8_1763_inst_req_0); -- 
    populateRxQueue_CP_2805_elements(18) <= populateRxQueue_CP_2805_elements(0);
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Sample/ra
      -- 
    ra_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u8_u8_1763_inst_ack_0, ack => populateRxQueue_CP_2805_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/Update/ca
      -- 
    ca_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u8_u8_1763_inst_ack_1, ack => populateRxQueue_CP_2805_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	25 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/$exit
      -- CP-element group 21: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/$exit
      -- CP-element group 21: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$exit
      -- CP-element group 21: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/$exit
      -- CP-element group 21: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_sources/AND_u8_u8_1763/SplitProtocol/$exit
      -- CP-element group 21: 	 branch_block_stmt_1752/merge_stmt_1753__entry___PhiReq/phi_stmt_1754/phi_stmt_1754_req
      -- 
    phi_stmt_1754_req_3087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1754_req_3087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(21), ack => phi_stmt_1754_req_0); -- 
    populateRxQueue_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_2805_elements(19) & populateRxQueue_CP_2805_elements(20);
      gj_populateRxQueue_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_2805_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	14 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Sample/ack
      -- 
    ack_3104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1785_1764_buf_ack_0, ack => populateRxQueue_CP_2805_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	14 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/Update/ack
      -- 
    ack_3109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1785_1764_buf_ack_1, ack => populateRxQueue_CP_2805_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_1752/loopback_PhiReq/$exit
      -- CP-element group 24: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/$exit
      -- CP-element group 24: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/$exit
      -- CP-element group 24: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_sources/Interlock/$exit
      -- CP-element group 24: 	 branch_block_stmt_1752/loopback_PhiReq/phi_stmt_1754/phi_stmt_1754_req
      -- 
    phi_stmt_1754_req_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1754_req_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(24), ack => phi_stmt_1754_req_1); -- 
    populateRxQueue_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_2805_elements(22) & populateRxQueue_CP_2805_elements(23);
      gj_populateRxQueue_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_2805_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  merge  transition  place  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	21 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1752/merge_stmt_1753_PhiReqMerge
      -- CP-element group 25: 	 branch_block_stmt_1752/merge_stmt_1753_PhiAck/$entry
      -- 
    populateRxQueue_CP_2805_elements(25) <= OrReduce(populateRxQueue_CP_2805_elements(21) & populateRxQueue_CP_2805_elements(24));
    -- CP-element group 26:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: 	3 
    -- CP-element group 26: 	5 
    -- CP-element group 26: 	6 
    -- CP-element group 26: 	7 
    -- CP-element group 26:  members (20) 
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Update/ccr
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Sample/crr
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Update/ccr
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1775_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/call_stmt_1773_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/$entry
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785__entry__
      -- CP-element group 26: 	 branch_block_stmt_1752/merge_stmt_1753__exit__
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1752/call_stmt_1773_to_assign_stmt_1785/AND_u8_u8_1784_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1752/merge_stmt_1753_PhiAck/$exit
      -- CP-element group 26: 	 branch_block_stmt_1752/merge_stmt_1753_PhiAck/phi_stmt_1754_ack
      -- 
    phi_stmt_1754_ack_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1754_ack_0, ack => populateRxQueue_CP_2805_elements(26)); -- 
    ccr_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(26), ack => call_stmt_1773_call_req_1); -- 
    crr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(26), ack => call_stmt_1773_call_req_0); -- 
    ccr_2848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(26), ack => call_stmt_1775_call_req_1); -- 
    cr_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(26), ack => AND_u8_u8_1784_inst_req_1); -- 
    rr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2805_elements(26), ack => AND_u8_u8_1784_inst_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_1758_wire : std_logic_vector(7 downto 0);
    signal ADD_u8_u8_1779_wire : std_logic_vector(7 downto 0);
    signal AND_u8_u8_1763_wire : std_logic_vector(7 downto 0);
    signal EQ_u1_u1_1798_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1791_wire : std_logic_vector(0 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756_wire : std_logic_vector(7 downto 0);
    signal RPIPE_S_NUMBER_OF_SERVERS_1759_wire : std_logic_vector(31 downto 0);
    signal RPIPE_S_NUMBER_OF_SERVERS_1780_wire : std_logic_vector(31 downto 0);
    signal R_RXQUEUE_1769_wire_constant : std_logic_vector(1 downto 0);
    signal SUB_u32_u32_1761_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1782_wire : std_logic_vector(31 downto 0);
    signal konst_1757_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1760_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1778_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1781_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1792_wire_constant : std_logic_vector(9 downto 0);
    signal konst_1797_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_1785 : std_logic_vector(7 downto 0);
    signal n_q_index_1785_1764_buffered : std_logic_vector(7 downto 0);
    signal push_status_1773 : std_logic_vector(0 downto 0);
    signal q_index_1754 : std_logic_vector(7 downto 0);
    signal status_1794 : std_logic_vector(0 downto 0);
    signal type_cast_1762_wire : std_logic_vector(7 downto 0);
    signal type_cast_1783_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_RXQUEUE_1769_wire_constant <= "10";
    konst_1757_wire_constant <= "00000001";
    konst_1760_wire_constant <= "00000000000000000000000000000001";
    konst_1778_wire_constant <= "00000001";
    konst_1781_wire_constant <= "00000000000000000000000000000001";
    konst_1792_wire_constant <= "0000100000";
    konst_1797_wire_constant <= "0";
    phi_stmt_1754: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= AND_u8_u8_1763_wire & n_q_index_1785_1764_buffered;
      req <= phi_stmt_1754_req_0 & phi_stmt_1754_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1754",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1754_ack_0,
          idata => idata,
          odata => q_index_1754,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1754
    n_q_index_1785_1764_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_1785_1764_buf_req_0;
      n_q_index_1785_1764_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_1785_1764_buf_req_1;
      n_q_index_1785_1764_buf_ack_1<= rack(0);
      n_q_index_1785_1764_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_1785_1764_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_1785,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_1785_1764_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1762_inst
    process(SUB_u32_u32_1761_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u32_u32_1761_wire(7 downto 0);
      type_cast_1762_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1783_inst
    process(SUB_u32_u32_1782_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u32_u32_1782_wire(7 downto 0);
      type_cast_1783_wire <= tmp_var; -- 
    end process;
    if_stmt_1789_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1791_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1789_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1789_branch_req_0,
          ack0 => if_stmt_1789_branch_ack_0,
          ack1 => if_stmt_1789_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1795_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_1798_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1795_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1795_branch_req_0,
          ack0 => if_stmt_1795_branch_ack_0,
          ack1 => if_stmt_1795_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u8_u8_1758_inst
    ADD_u8_u8_1758_wire <= std_logic_vector(unsigned(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756_wire) + unsigned(konst_1757_wire_constant));
    -- flow through binary operator ADD_u8_u8_1779_inst
    ADD_u8_u8_1779_wire <= std_logic_vector(unsigned(q_index_1754) + unsigned(konst_1778_wire_constant));
    -- shared split operator group (2) : AND_u8_u8_1763_inst 
    ApIntAnd_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u8_u8_1758_wire & type_cast_1762_wire;
      AND_u8_u8_1763_wire <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u8_u8_1763_inst_req_0;
      AND_u8_u8_1763_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u8_u8_1763_inst_req_1;
      AND_u8_u8_1763_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : AND_u8_u8_1784_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u8_u8_1779_wire & type_cast_1783_wire;
      n_q_index_1785 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u8_u8_1784_inst_req_0;
      AND_u8_u8_1784_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u8_u8_1784_inst_req_1;
      AND_u8_u8_1784_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- flow through binary operator EQ_u1_u1_1798_inst
    process(status_1794) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_1794, konst_1797_wire_constant, tmp_var);
      EQ_u1_u1_1798_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1791_inst
    process(push_status_1773) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_1773, tmp_var);
      NOT_u1_u1_1791_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator SUB_u32_u32_1761_inst
    SUB_u32_u32_1761_wire <= std_logic_vector(unsigned(RPIPE_S_NUMBER_OF_SERVERS_1759_wire) - unsigned(konst_1760_wire_constant));
    -- flow through binary operator SUB_u32_u32_1782_inst
    SUB_u32_u32_1782_wire <= std_logic_vector(unsigned(RPIPE_S_NUMBER_OF_SERVERS_1780_wire) - unsigned(konst_1781_wire_constant));
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1756_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- read from input-signal S_NUMBER_OF_SERVERS
    RPIPE_S_NUMBER_OF_SERVERS_1759_wire <= S_NUMBER_OF_SERVERS;
    RPIPE_S_NUMBER_OF_SERVERS_1780_wire <= S_NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1802_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_1754;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1773_call 
    pushIntoQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(81 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1773_call_req_0;
      call_stmt_1773_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1773_call_req_1;
      call_stmt_1773_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_0_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_RXQUEUE_1769_wire_constant & q_index_1754 & rx_buffer_pointer_buffer;
      push_status_1773 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 82,
        owidth => 82,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(81 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1775_call 
    incrementNumberOfPacketsReceived_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1775_call_req_0;
      call_stmt_1775_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1775_call_req_1;
      call_stmt_1775_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not push_status_1773(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      incrementNumberOfPacketsReceived_call_group_1_gI: SplitGuardInterface generic map(name => "incrementNumberOfPacketsReceived_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => incrementNumberOfPacketsReceived_call_reqs(0),
          ackR => incrementNumberOfPacketsReceived_call_acks(0),
          tagR => incrementNumberOfPacketsReceived_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => incrementNumberOfPacketsReceived_return_acks(0), -- cross-over
          ackL => incrementNumberOfPacketsReceived_return_reqs(0), -- cross-over
          tagL => incrementNumberOfPacketsReceived_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    operator_delay_time_4570_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_1794_call_req_0;
      call_stmt_1794_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_1794_call_req_1;
      call_stmt_1794_call_ack_1<= update_ack(0);
      call_stmt_1794_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_1792_wire_constant,
        delay_done => status_1794,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    queue_type : in  std_logic_vector(1 downto 0);
    server_id : in  std_logic_vector(7 downto 0);
    q_w_data : in  std_logic_vector(63 downto 0);
    status : out  std_logic_vector(0 downto 0);
    QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
    QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
    QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
    getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
    getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
    getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
    getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
    accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
    accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(71 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
    setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(71 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
    getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
    getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
    getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
    getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(71 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(167 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 82)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal queue_type_buffer :  std_logic_vector(1 downto 0);
  signal queue_type_update_enable: Boolean;
  signal server_id_buffer :  std_logic_vector(7 downto 0);
  signal server_id_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(63 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_2429_start: Boolean;
  signal pushIntoQueue_CP_2429_symbol: Boolean;
  -- volatile/operator module components. 
  component getQueuePointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLockPointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock_address_pointer : in  std_logic_vector(63 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_data : out  std_logic_vector(135 downto 0);
      accessMemoryLdStub_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryLdStub_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
      accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      queue_length : out  std_logic_vector(31 downto 0);
      accessQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueLength_call_data : out  std_logic_vector(104 downto 0);
      accessQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueLength_return_data : in   std_logic_vector(31 downto 0);
      accessQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueBufPointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
      accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock_address_pointer : in  std_logic_vector(63 downto 0);
      accessMemoryByte_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByte_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByte_call_data : out  std_logic_vector(144 downto 0);
      accessMemoryByte_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryByte_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByte_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByte_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByte_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      buf_base_address : in  std_logic_vector(63 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(63 downto 0);
      accessQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_call_data : out  std_logic_vector(168 downto 0);
      accessQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_return_data : in   std_logic_vector(63 downto 0);
      accessQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1583_call_ack_0 : boolean;
  signal call_stmt_1591_call_req_0 : boolean;
  signal call_stmt_1591_call_ack_0 : boolean;
  signal call_stmt_1583_call_req_1 : boolean;
  signal call_stmt_1583_call_ack_1 : boolean;
  signal call_stmt_1583_call_req_0 : boolean;
  signal call_stmt_1591_call_req_1 : boolean;
  signal call_stmt_1591_call_ack_1 : boolean;
  signal call_stmt_1601_call_req_0 : boolean;
  signal call_stmt_1601_call_ack_0 : boolean;
  signal call_stmt_1601_call_req_1 : boolean;
  signal call_stmt_1601_call_ack_1 : boolean;
  signal call_stmt_1606_call_req_0 : boolean;
  signal call_stmt_1606_call_ack_0 : boolean;
  signal call_stmt_1606_call_req_1 : boolean;
  signal call_stmt_1606_call_ack_1 : boolean;
  signal call_stmt_1612_call_req_0 : boolean;
  signal call_stmt_1612_call_ack_0 : boolean;
  signal call_stmt_1612_call_req_1 : boolean;
  signal call_stmt_1612_call_ack_1 : boolean;
  signal call_stmt_1616_call_req_0 : boolean;
  signal call_stmt_1616_call_ack_0 : boolean;
  signal call_stmt_1616_call_req_1 : boolean;
  signal call_stmt_1616_call_ack_1 : boolean;
  signal call_stmt_1620_call_req_0 : boolean;
  signal call_stmt_1620_call_ack_0 : boolean;
  signal call_stmt_1620_call_req_1 : boolean;
  signal call_stmt_1620_call_ack_1 : boolean;
  signal call_stmt_1645_call_req_0 : boolean;
  signal call_stmt_1645_call_ack_0 : boolean;
  signal call_stmt_1645_call_req_1 : boolean;
  signal call_stmt_1645_call_ack_1 : boolean;
  signal call_stmt_1651_call_req_0 : boolean;
  signal call_stmt_1651_call_ack_0 : boolean;
  signal call_stmt_1651_call_req_1 : boolean;
  signal call_stmt_1651_call_ack_1 : boolean;
  signal call_stmt_1657_call_req_0 : boolean;
  signal call_stmt_1657_call_ack_0 : boolean;
  signal call_stmt_1657_call_req_1 : boolean;
  signal call_stmt_1657_call_ack_1 : boolean;
  signal call_stmt_1665_call_req_0 : boolean;
  signal call_stmt_1665_call_ack_0 : boolean;
  signal call_stmt_1665_call_req_1 : boolean;
  signal call_stmt_1665_call_ack_1 : boolean;
  signal CONCAT_u16_u32_1682_inst_req_0 : boolean;
  signal CONCAT_u16_u32_1682_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_1682_inst_req_1 : boolean;
  signal CONCAT_u16_u32_1682_inst_ack_1 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_req_0 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_ack_0 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_req_1 : boolean;
  signal WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_ack_1 : boolean;
  signal call_stmt_1688_call_req_0 : boolean;
  signal call_stmt_1688_call_ack_0 : boolean;
  signal call_stmt_1688_call_req_1 : boolean;
  signal call_stmt_1688_call_ack_1 : boolean;
  signal W_status_1689_inst_req_0 : boolean;
  signal W_status_1689_inst_ack_0 : boolean;
  signal W_status_1689_inst_req_1 : boolean;
  signal W_status_1689_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 82) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(9 downto 8) <= queue_type;
  queue_type_buffer <= in_buffer_data_out(9 downto 8);
  in_buffer_data_in(17 downto 10) <= server_id;
  server_id_buffer <= in_buffer_data_out(17 downto 10);
  in_buffer_data_in(81 downto 18) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(81 downto 18);
  in_buffer_data_in(tag_length + 81 downto 82) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 81 downto 82);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_2429_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_2429_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_2429_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_2429_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_2429: Block -- control-path 
    signal pushIntoQueue_CP_2429_elements: BooleanArray(41 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_2429_elements(0) <= pushIntoQueue_CP_2429_start;
    pushIntoQueue_CP_2429_symbol <= pushIntoQueue_CP_2429_elements(41);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/$entry
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Update/$entry
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Update/$entry
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Update/ccr
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_update_start_
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_update_start_
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_sample_start_
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Sample/crr
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Update/ccr
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_update_start_
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Update/$entry
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Update/ccr
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_update_start_
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Update/$entry
      -- CP-element group 0: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Update/ccr
      -- 
    crr_2442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(0), ack => call_stmt_1583_call_req_0); -- 
    ccr_2447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(0), ack => call_stmt_1583_call_req_1); -- 
    ccr_2461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(0), ack => call_stmt_1591_call_req_1); -- 
    ccr_2475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(0), ack => call_stmt_1601_call_req_1); -- 
    ccr_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(0), ack => call_stmt_1606_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Sample/cra
      -- CP-element group 1: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_sample_completed_
      -- CP-element group 1: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Sample/$exit
      -- 
    cra_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1583_call_ack_0, ack => pushIntoQueue_CP_2429_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	11 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Sample/crr
      -- CP-element group 2: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Update/$exit
      -- CP-element group 2: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_Update/cca
      -- CP-element group 2: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_update_completed_
      -- CP-element group 2: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_sample_start_
      -- 
    cca_2448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1583_call_ack_1, ack => pushIntoQueue_CP_2429_elements(2)); -- 
    crr_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(2), ack => call_stmt_1591_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Sample/cra
      -- CP-element group 3: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_sample_completed_
      -- CP-element group 3: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Sample/$exit
      -- 
    cra_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1591_call_ack_0, ack => pushIntoQueue_CP_2429_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	8 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Update/$exit
      -- CP-element group 4: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_update_completed_
      -- CP-element group 4: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1591_Update/cca
      -- 
    cca_2462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1591_call_ack_1, ack => pushIntoQueue_CP_2429_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	11 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_sample_start_
      -- CP-element group 5: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Sample/$entry
      -- CP-element group 5: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Sample/crr
      -- 
    crr_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(5), ack => call_stmt_1601_call_req_0); -- 
    pushIntoQueue_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "pushIntoQueue_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(4) & pushIntoQueue_CP_2429_elements(11);
      gj_pushIntoQueue_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_sample_completed_
      -- CP-element group 6: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Sample/$exit
      -- CP-element group 6: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Sample/cra
      -- 
    cra_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1601_call_ack_0, ack => pushIntoQueue_CP_2429_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_update_completed_
      -- CP-element group 7: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Update/$exit
      -- CP-element group 7: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1601_Update/cca
      -- 
    cca_2476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1601_call_ack_1, ack => pushIntoQueue_CP_2429_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_sample_start_
      -- CP-element group 8: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Sample/crr
      -- 
    crr_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(8), ack => call_stmt_1606_call_req_0); -- 
    pushIntoQueue_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "pushIntoQueue_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(4) & pushIntoQueue_CP_2429_elements(7);
      gj_pushIntoQueue_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_sample_completed_
      -- CP-element group 9: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Sample/$exit
      -- CP-element group 9: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Sample/cra
      -- 
    cra_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1606_call_ack_0, ack => pushIntoQueue_CP_2429_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	26 
    -- CP-element group 10: 	29 
    -- CP-element group 10: 	32 
    -- CP-element group 10:  members (32) 
      -- CP-element group 10: 	 call_stmt_1583_to_call_stmt_1606/$exit
      -- CP-element group 10: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_update_completed_
      -- CP-element group 10: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Update/$exit
      -- CP-element group 10: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1606_Update/cca
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_sample_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Sample/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Sample/crr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Update/ccr
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_update_start_
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Update/$entry
      -- CP-element group 10: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Update/cr
      -- 
    cca_2490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1606_call_ack_1, ack => pushIntoQueue_CP_2429_elements(10)); -- 
    crr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1612_call_req_0); -- 
    ccr_2507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1612_call_req_1); -- 
    ccr_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1616_call_req_1); -- 
    ccr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1620_call_req_1); -- 
    ccr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1645_call_req_1); -- 
    ccr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1651_call_req_1); -- 
    ccr_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1657_call_req_1); -- 
    ccr_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => call_stmt_1665_call_req_1); -- 
    cr_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(10), ack => CONCAT_u16_u32_1682_inst_req_1); -- 
    -- CP-element group 11:  transition  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	5 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 call_stmt_1583_to_call_stmt_1606/call_stmt_1583_call_stmt_1601_delay
      -- 
    -- Element group pushIntoQueue_CP_2429_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => pushIntoQueue_CP_2429_elements(2), ack => pushIntoQueue_CP_2429_elements(11), clk => clk, reset =>reset);
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_sample_completed_
      -- CP-element group 12: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Sample/$exit
      -- CP-element group 12: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Sample/cra
      -- 
    cra_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1612_call_ack_0, ack => pushIntoQueue_CP_2429_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	21 
    -- CP-element group 13: 	24 
    -- CP-element group 13: 	30 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_update_completed_
      -- CP-element group 13: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Update/$exit
      -- CP-element group 13: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1612_Update/cca
      -- CP-element group 13: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_sample_start_
      -- CP-element group 13: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Sample/$entry
      -- CP-element group 13: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Sample/crr
      -- 
    cca_2508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1612_call_ack_1, ack => pushIntoQueue_CP_2429_elements(13)); -- 
    crr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(13), ack => call_stmt_1616_call_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_sample_completed_
      -- CP-element group 14: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Sample/$exit
      -- CP-element group 14: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Sample/cra
      -- 
    cra_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1616_call_ack_0, ack => pushIntoQueue_CP_2429_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	33 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_update_completed_
      -- CP-element group 15: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Update/$exit
      -- CP-element group 15: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1616_Update/cca
      -- CP-element group 15: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_sample_start_
      -- CP-element group 15: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Sample/$entry
      -- CP-element group 15: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Sample/crr
      -- 
    cca_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1616_call_ack_1, ack => pushIntoQueue_CP_2429_elements(15)); -- 
    crr_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(15), ack => call_stmt_1620_call_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_sample_completed_
      -- CP-element group 16: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Sample/$exit
      -- CP-element group 16: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Sample/cra
      -- 
    cra_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1620_call_ack_0, ack => pushIntoQueue_CP_2429_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	27 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	33 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_update_completed_
      -- CP-element group 17: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Update/$exit
      -- CP-element group 17: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1620_Update/cca
      -- 
    cca_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1620_call_ack_1, ack => pushIntoQueue_CP_2429_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_sample_start_
      -- CP-element group 18: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Sample/$entry
      -- CP-element group 18: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Sample/crr
      -- 
    crr_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(18), ack => call_stmt_1645_call_req_0); -- 
    pushIntoQueue_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(15) & pushIntoQueue_CP_2429_elements(17);
      gj_pushIntoQueue_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_sample_completed_
      -- CP-element group 19: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Sample/$exit
      -- CP-element group 19: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Sample/cra
      -- 
    cra_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1645_call_ack_0, ack => pushIntoQueue_CP_2429_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_update_completed_
      -- CP-element group 20: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Update/$exit
      -- CP-element group 20: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1645_Update/cca
      -- 
    cca_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1645_call_ack_1, ack => pushIntoQueue_CP_2429_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	13 
    -- CP-element group 21: 	15 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_sample_start_
      -- CP-element group 21: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Sample/$entry
      -- CP-element group 21: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Sample/crr
      -- 
    crr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(21), ack => call_stmt_1651_call_req_0); -- 
    pushIntoQueue_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(13) & pushIntoQueue_CP_2429_elements(15) & pushIntoQueue_CP_2429_elements(17) & pushIntoQueue_CP_2429_elements(20);
      gj_pushIntoQueue_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_sample_completed_
      -- CP-element group 22: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Sample/$exit
      -- CP-element group 22: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Sample/cra
      -- 
    cra_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1651_call_ack_0, ack => pushIntoQueue_CP_2429_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_update_completed_
      -- CP-element group 23: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Update/$exit
      -- CP-element group 23: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1651_Update/cca
      -- 
    cca_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1651_call_ack_1, ack => pushIntoQueue_CP_2429_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	13 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	17 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_sample_start_
      -- CP-element group 24: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Sample/$entry
      -- CP-element group 24: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Sample/crr
      -- 
    crr_2572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(24), ack => call_stmt_1657_call_req_0); -- 
    pushIntoQueue_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(13) & pushIntoQueue_CP_2429_elements(15) & pushIntoQueue_CP_2429_elements(17) & pushIntoQueue_CP_2429_elements(23);
      gj_pushIntoQueue_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_sample_completed_
      -- CP-element group 25: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Sample/$exit
      -- CP-element group 25: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Sample/cra
      -- 
    cra_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1657_call_ack_0, ack => pushIntoQueue_CP_2429_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	10 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_update_completed_
      -- CP-element group 26: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Update/$exit
      -- CP-element group 26: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1657_Update/cca
      -- 
    cca_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1657_call_ack_1, ack => pushIntoQueue_CP_2429_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: 	17 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_sample_start_
      -- CP-element group 27: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Sample/$entry
      -- CP-element group 27: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Sample/crr
      -- 
    crr_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(27), ack => call_stmt_1665_call_req_0); -- 
    pushIntoQueue_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(15) & pushIntoQueue_CP_2429_elements(17) & pushIntoQueue_CP_2429_elements(26);
      gj_pushIntoQueue_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_sample_completed_
      -- CP-element group 28: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Sample/$exit
      -- CP-element group 28: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Sample/cra
      -- 
    cra_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1665_call_ack_0, ack => pushIntoQueue_CP_2429_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	10 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	36 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_update_completed_
      -- CP-element group 29: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Update/$exit
      -- CP-element group 29: 	 call_stmt_1612_to_assign_stmt_1683/call_stmt_1665_Update/cca
      -- 
    cca_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1665_call_ack_1, ack => pushIntoQueue_CP_2429_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	13 
    -- CP-element group 30: 	15 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_sample_start_
      -- CP-element group 30: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Sample/$entry
      -- CP-element group 30: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Sample/rr
      -- 
    rr_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(30), ack => CONCAT_u16_u32_1682_inst_req_0); -- 
    pushIntoQueue_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(13) & pushIntoQueue_CP_2429_elements(15) & pushIntoQueue_CP_2429_elements(17);
      gj_pushIntoQueue_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_sample_completed_
      -- CP-element group 31: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Sample/$exit
      -- CP-element group 31: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Sample/ra
      -- 
    ra_2601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1682_inst_ack_0, ack => pushIntoQueue_CP_2429_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	10 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_update_completed_
      -- CP-element group 32: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Update/$exit
      -- CP-element group 32: 	 call_stmt_1612_to_assign_stmt_1683/CONCAT_u16_u32_1682_Update/ca
      -- 
    ca_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_1682_inst_ack_1, ack => pushIntoQueue_CP_2429_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: 	17 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_sample_start_
      -- CP-element group 33: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Sample/$entry
      -- CP-element group 33: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Sample/req
      -- 
    req_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(33), ack => WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_req_0); -- 
    pushIntoQueue_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(15) & pushIntoQueue_CP_2429_elements(17) & pushIntoQueue_CP_2429_elements(32);
      gj_pushIntoQueue_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_sample_completed_
      -- CP-element group 34: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_update_start_
      -- CP-element group 34: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Sample/$exit
      -- CP-element group 34: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Sample/ack
      -- CP-element group 34: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Update/$entry
      -- CP-element group 34: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Update/req
      -- 
    ack_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_ack_0, ack => pushIntoQueue_CP_2429_elements(34)); -- 
    req_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(34), ack => WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_update_completed_
      -- CP-element group 35: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Update/$exit
      -- CP-element group 35: 	 call_stmt_1612_to_assign_stmt_1683/WPIPE_QUEUE_MONITOR_SIGNAL_1667_Update/ack
      -- 
    ack_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_ack_1, ack => pushIntoQueue_CP_2429_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	29 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36: 	39 
    -- CP-element group 36: 	40 
    -- CP-element group 36:  members (14) 
      -- CP-element group 36: 	 call_stmt_1612_to_assign_stmt_1683/$exit
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/$entry
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_sample_start_
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_update_start_
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Sample/$entry
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Sample/crr
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Update/$entry
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Update/ccr
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_sample_start_
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_update_start_
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Sample/$entry
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Sample/req
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Update/$entry
      -- CP-element group 36: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Update/req
      -- 
    crr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(36), ack => call_stmt_1688_call_req_0); -- 
    ccr_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(36), ack => call_stmt_1688_call_req_1); -- 
    req_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(36), ack => W_status_1689_inst_req_0); -- 
    req_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_2429_elements(36), ack => W_status_1689_inst_req_1); -- 
    pushIntoQueue_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(29) & pushIntoQueue_CP_2429_elements(35);
      gj_pushIntoQueue_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_sample_completed_
      -- CP-element group 37: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Sample/$exit
      -- CP-element group 37: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Sample/cra
      -- 
    cra_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1688_call_ack_0, ack => pushIntoQueue_CP_2429_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_update_completed_
      -- CP-element group 38: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Update/$exit
      -- CP-element group 38: 	 call_stmt_1688_to_assign_stmt_1691/call_stmt_1688_Update/cca
      -- 
    cca_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1688_call_ack_1, ack => pushIntoQueue_CP_2429_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	36 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_sample_completed_
      -- CP-element group 39: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Sample/$exit
      -- CP-element group 39: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Sample/ack
      -- 
    ack_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1689_inst_ack_0, ack => pushIntoQueue_CP_2429_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	36 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_update_completed_
      -- CP-element group 40: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Update/$exit
      -- CP-element group 40: 	 call_stmt_1688_to_assign_stmt_1691/assign_stmt_1691_Update/ack
      -- 
    ack_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1689_inst_ack_1, ack => pushIntoQueue_CP_2429_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 $exit
      -- CP-element group 41: 	 call_stmt_1688_to_assign_stmt_1691/$exit
      -- 
    pushIntoQueue_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_2429_elements(38) & pushIntoQueue_CP_2429_elements(40);
      gj_pushIntoQueue_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_2429_elements(41), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1633_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1664_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1674_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1682_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u4_u8_1671_wire : std_logic_vector(7 downto 0);
    signal CONCAT_u8_u16_1676_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_1681_wire : std_logic_vector(15 downto 0);
    signal R_PUSHQ_1670_wire_constant : std_logic_vector(3 downto 0);
    signal R_READMEM_1585_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u32_u32_1625_wire : std_logic_vector(31 downto 0);
    signal konst_1587_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1594_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1624_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1630_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1632_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1673_wire_constant : std_logic_vector(31 downto 0);
    signal lock_n_1596 : std_logic_vector(0 downto 0);
    signal m_ok_1606 : std_logic_vector(0 downto 0);
    signal misc_1591 : std_logic_vector(31 downto 0);
    signal next_wi_1635 : std_logic_vector(31 downto 0);
    signal q_base_address_1583 : std_logic_vector(63 downto 0);
    signal q_buf_address_1645 : std_logic_vector(63 downto 0);
    signal q_full_1640 : std_logic_vector(0 downto 0);
    signal q_lock_address_1601 : std_logic_vector(63 downto 0);
    signal queue_length_1616 : std_logic_vector(31 downto 0);
    signal read_index_1612 : std_logic_vector(31 downto 0);
    signal round_off_1627 : std_logic_vector(0 downto 0);
    signal total_msgs_1620 : std_logic_vector(31 downto 0);
    signal type_cast_1589_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1663_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1669_wire : std_logic_vector(3 downto 0);
    signal type_cast_1675_wire : std_logic_vector(7 downto 0);
    signal type_cast_1678_wire : std_logic_vector(7 downto 0);
    signal type_cast_1680_wire : std_logic_vector(7 downto 0);
    signal write_index_1612 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_PUSHQ_1670_wire_constant <= "0010";
    R_READMEM_1585_wire_constant <= "1";
    konst_1587_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011100";
    konst_1594_wire_constant <= "00000000000000000000000000000000";
    konst_1624_wire_constant <= "00000000000000000000000000000001";
    konst_1630_wire_constant <= "00000000000000000000000000000000";
    konst_1632_wire_constant <= "00000000000000000000000000000001";
    konst_1673_wire_constant <= "00000000000000000000000000000001";
    type_cast_1589_wire_constant <= "00000000000000000000000000000000";
    type_cast_1663_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_1634_inst
    next_wi_1635 <= konst_1630_wire_constant when (round_off_1627(0) /=  '0') else ADD_u32_u32_1633_wire;
    W_status_1689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_1689_inst_req_0;
      W_status_1689_inst_ack_0<= wack(0);
      rreq(0) <= W_status_1689_inst_req_1;
      W_status_1689_inst_ack_1<= rack(0);
      W_status_1689_inst : InterlockBuffer generic map ( -- 
        name => "W_status_1689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_full_1640,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1669_inst
    process(queue_type_buffer) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := queue_type_buffer(1 downto 0);
      type_cast_1669_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1675_inst
    process(ADD_u32_u32_1674_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ADD_u32_u32_1674_wire(7 downto 0);
      type_cast_1675_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1678_inst
    process(next_wi_1635) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := next_wi_1635(7 downto 0);
      type_cast_1678_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1680_inst
    process(read_index_1612) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := read_index_1612(7 downto 0);
      type_cast_1680_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator ADD_u32_u32_1633_inst
    ADD_u32_u32_1633_wire <= std_logic_vector(unsigned(write_index_1612) + unsigned(konst_1632_wire_constant));
    -- flow through binary operator ADD_u32_u32_1664_inst
    ADD_u32_u32_1664_wire <= std_logic_vector(unsigned(total_msgs_1620) + unsigned(type_cast_1663_wire_constant));
    -- flow through binary operator ADD_u32_u32_1674_inst
    ADD_u32_u32_1674_wire <= std_logic_vector(unsigned(total_msgs_1620) + unsigned(konst_1673_wire_constant));
    -- flow through binary operator BITSEL_u32_u1_1595_inst
    process(misc_1591) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(misc_1591, konst_1594_wire_constant, tmp_var);
      lock_n_1596 <= tmp_var; --
    end process;
    -- shared split operator group (4) : CONCAT_u16_u32_1682_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_1676_wire & CONCAT_u8_u16_1681_wire;
      CONCAT_u16_u32_1682_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  not q_full_1640(0);
      reqL_unguarded(0) <= CONCAT_u16_u32_1682_inst_req_0;
      CONCAT_u16_u32_1682_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_1682_inst_req_1;
      CONCAT_u16_u32_1682_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- flow through binary operator CONCAT_u4_u8_1671_inst
    process(type_cast_1669_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1669_wire, R_PUSHQ_1670_wire_constant, tmp_var);
      CONCAT_u4_u8_1671_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_1676_inst
    process(CONCAT_u4_u8_1671_wire, type_cast_1675_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u8_1671_wire, type_cast_1675_wire, tmp_var);
      CONCAT_u8_u16_1676_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u8_u16_1681_inst
    process(type_cast_1678_wire, type_cast_1680_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1678_wire, type_cast_1680_wire, tmp_var);
      CONCAT_u8_u16_1681_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_1626_inst
    process(write_index_1612, SUB_u32_u32_1625_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_1612, SUB_u32_u32_1625_wire, tmp_var);
      round_off_1627 <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_1639_inst
    process(total_msgs_1620, queue_length_1616) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(total_msgs_1620, queue_length_1616, tmp_var);
      q_full_1640 <= tmp_var; --
    end process;
    -- flow through binary operator SUB_u32_u32_1625_inst
    SUB_u32_u32_1625_wire <= std_logic_vector(unsigned(queue_length_1616) - unsigned(konst_1624_wire_constant));
    -- shared outport operator group (0) : WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_req_0;
      WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_req_1;
      WPIPE_QUEUE_MONITOR_SIGNAL_1667_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not q_full_1640(0);
      data_in <= CONCAT_u16_u32_1682_wire;
      QUEUE_MONITOR_SIGNAL_write_0_gI: SplitGuardInterface generic map(name => "QUEUE_MONITOR_SIGNAL_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      QUEUE_MONITOR_SIGNAL_write_0: OutputPortRevised -- 
        generic map ( name => "QUEUE_MONITOR_SIGNAL", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => QUEUE_MONITOR_SIGNAL_pipe_write_req(0),
          oack => QUEUE_MONITOR_SIGNAL_pipe_write_ack(0),
          odata => QUEUE_MONITOR_SIGNAL_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1583_call 
    getQueuePointer_call_group_0: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1583_call_req_0;
      call_stmt_1583_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1583_call_req_1;
      call_stmt_1583_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointer_call_group_0_gI: SplitGuardInterface generic map(name => "getQueuePointer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= queue_type_buffer & server_id_buffer;
      q_base_address_1583 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 10,
        owidth => 10,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointer_call_reqs(0),
          ackR => getQueuePointer_call_acks(0),
          dataR => getQueuePointer_call_data(9 downto 0),
          tagR => getQueuePointer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointer_return_acks(0), -- cross-over
          ackL => getQueuePointer_return_reqs(0), -- cross-over
          dataL => getQueuePointer_return_data(63 downto 0),
          tagL => getQueuePointer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1591_call 
    accessMemoryWord_call_group_1: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1591_call_req_0;
      call_stmt_1591_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1591_call_req_1;
      call_stmt_1591_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryWord_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryWord_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_1585_wire_constant & q_base_address_1583 & konst_1587_wire_constant & type_cast_1589_wire_constant;
      misc_1591 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryWord_call_reqs(0),
          ackR => accessMemoryWord_call_acks(0),
          dataR => accessMemoryWord_call_data(168 downto 0),
          tagR => accessMemoryWord_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryWord_return_acks(0), -- cross-over
          ackL => accessMemoryWord_return_reqs(0), -- cross-over
          dataL => accessMemoryWord_return_data(31 downto 0),
          tagL => accessMemoryWord_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1601_call 
    getQueueLockPointer_call_group_2: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1601_call_req_0;
      call_stmt_1601_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1601_call_req_1;
      call_stmt_1601_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not lock_n_1596(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLockPointer_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueLockPointer_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= queue_type_buffer & server_id_buffer;
      q_lock_address_1601 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 10,
        owidth => 10,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLockPointer_call_reqs(0),
          ackR => getQueueLockPointer_call_acks(0),
          dataR => getQueueLockPointer_call_data(9 downto 0),
          tagR => getQueueLockPointer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLockPointer_return_acks(0), -- cross-over
          ackL => getQueueLockPointer_return_reqs(0), -- cross-over
          dataL => getQueueLockPointer_return_data(63 downto 0),
          tagL => getQueueLockPointer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1606_call 
    acquireLock_call_group_3: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1606_call_req_0;
      call_stmt_1606_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1606_call_req_1;
      call_stmt_1606_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not lock_n_1596(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_3_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_lock_address_1601;
      m_ok_1606 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(71 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1612_call 
    getQueuePointers_call_group_4: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1612_call_req_0;
      call_stmt_1612_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1612_call_req_1;
      call_stmt_1612_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_4_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1583;
      write_index_1612 <= data_out(63 downto 32);
      read_index_1612 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(71 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1616_call 
    getQueueLength_call_group_5: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1616_call_req_0;
      call_stmt_1616_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1616_call_req_1;
      call_stmt_1616_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_5_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1583;
      queue_length_1616 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(71 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1620_call 
    getTotalMessages_call_group_6: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1620_call_req_0;
      call_stmt_1620_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1620_call_req_1;
      call_stmt_1620_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_6_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1583;
      total_msgs_1620 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(71 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1645_call 
    getQueueBufPointer_call_group_7: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1645_call_req_0;
      call_stmt_1645_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1645_call_req_1;
      call_stmt_1645_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1640(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueBufPointer_call_group_7_gI: SplitGuardInterface generic map(name => "getQueueBufPointer_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= queue_type_buffer & server_id_buffer;
      q_buf_address_1645 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 10,
        owidth => 10,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueBufPointer_call_reqs(0),
          ackR => getQueueBufPointer_call_acks(0),
          dataR => getQueueBufPointer_call_data(9 downto 0),
          tagR => getQueueBufPointer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueBufPointer_return_acks(0), -- cross-over
          ackL => getQueueBufPointer_return_reqs(0), -- cross-over
          dataL => getQueueBufPointer_return_data(63 downto 0),
          tagL => getQueueBufPointer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_1651_call 
    setQueueElement_call_group_8: Block -- 
      signal data_in: std_logic_vector(167 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1651_call_req_0;
      call_stmt_1651_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1651_call_req_1;
      call_stmt_1651_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1640(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_8_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_buf_address_1645 & write_index_1612 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 168,
        owidth => 168,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(167 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- shared call operator group (9) : call_stmt_1657_call 
    setQueuePointers_call_group_9: Block -- 
      signal data_in: std_logic_vector(135 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1657_call_req_0;
      call_stmt_1657_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1657_call_req_1;
      call_stmt_1657_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1640(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_9_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1583 & next_wi_1635 & read_index_1612;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 136,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(135 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 9
    -- shared call operator group (10) : call_stmt_1665_call 
    setTotalMessages_call_group_10: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1665_call_req_0;
      call_stmt_1665_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1665_call_req_1;
      call_stmt_1665_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1640(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setTotalMessages_call_group_10_gI: SplitGuardInterface generic map(name => "setTotalMessages_call_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_base_address_1583 & ADD_u32_u32_1664_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setTotalMessages_call_reqs(0),
          ackR => setTotalMessages_call_acks(0),
          dataR => setTotalMessages_call_data(103 downto 0),
          tagR => setTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setTotalMessages_return_acks(0), -- cross-over
          ackL => setTotalMessages_return_reqs(0), -- cross-over
          tagL => setTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 10
    -- shared call operator group (11) : call_stmt_1688_call 
    releaseLock_call_group_11: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1688_call_req_0;
      call_stmt_1688_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1688_call_req_1;
      call_stmt_1688_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not lock_n_1596(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_11_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & q_lock_address_1601;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(71 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 11
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity releaseLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    lock_address_pointer : in  std_logic_vector(63 downto 0);
    accessMemoryByte_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryByte_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryByte_call_data : out  std_logic_vector(144 downto 0);
    accessMemoryByte_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMemoryByte_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryByte_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryByte_return_data : in   std_logic_vector(7 downto 0);
    accessMemoryByte_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseLock;
architecture releaseLock_arch of releaseLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal lock_address_pointer_buffer :  std_logic_vector(63 downto 0);
  signal lock_address_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal releaseLock_CP_1649_start: Boolean;
  signal releaseLock_CP_1649_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryByte is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      byte_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wbyte : in  std_logic_vector(7 downto 0);
      rbyte : out  std_logic_vector(7 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1197_call_req_0 : boolean;
  signal call_stmt_1197_call_ack_0 : boolean;
  signal call_stmt_1197_call_req_1 : boolean;
  signal call_stmt_1197_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= lock_address_pointer;
  lock_address_pointer_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseLock_CP_1649_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_1649_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseLock_CP_1649_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_1649_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseLock_CP_1649: Block -- control-path 
    signal releaseLock_CP_1649_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    releaseLock_CP_1649_elements(0) <= releaseLock_CP_1649_start;
    releaseLock_CP_1649_symbol <= releaseLock_CP_1649_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1197/$entry
      -- CP-element group 0: 	 call_stmt_1197/call_stmt_1197_sample_start_
      -- CP-element group 0: 	 call_stmt_1197/call_stmt_1197_update_start_
      -- CP-element group 0: 	 call_stmt_1197/call_stmt_1197_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1197/call_stmt_1197_Sample/crr
      -- CP-element group 0: 	 call_stmt_1197/call_stmt_1197_Update/$entry
      -- CP-element group 0: 	 call_stmt_1197/call_stmt_1197_Update/ccr
      -- 
    ccr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_1649_elements(0), ack => call_stmt_1197_call_req_1); -- 
    crr_1662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_1649_elements(0), ack => call_stmt_1197_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1197/call_stmt_1197_sample_completed_
      -- CP-element group 1: 	 call_stmt_1197/call_stmt_1197_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1197/call_stmt_1197_Sample/cra
      -- 
    cra_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1197_call_ack_0, ack => releaseLock_CP_1649_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1197/$exit
      -- CP-element group 2: 	 call_stmt_1197/call_stmt_1197_update_completed_
      -- CP-element group 2: 	 call_stmt_1197/call_stmt_1197_Update/$exit
      -- CP-element group 2: 	 call_stmt_1197/call_stmt_1197_Update/cca
      -- 
    cca_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1197_call_ack_1, ack => releaseLock_CP_1649_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_WRITEMEM_1192_wire_constant : std_logic_vector(0 downto 0);
    signal ignore_1197 : std_logic_vector(7 downto 0);
    signal konst_1194_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1195_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_WRITEMEM_1192_wire_constant <= "0";
    konst_1194_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_1195_wire_constant <= "00000000";
    -- shared call operator group (0) : call_stmt_1197_call 
    accessMemoryByte_call_group_0: Block -- 
      signal data_in: std_logic_vector(144 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1197_call_req_0;
      call_stmt_1197_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1197_call_req_1;
      call_stmt_1197_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryByte_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryByte_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_WRITEMEM_1192_wire_constant & lock_address_pointer_buffer & konst_1194_wire_constant & konst_1195_wire_constant;
      ignore_1197 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 145,
        owidth => 145,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryByte_call_reqs(0),
          ackR => accessMemoryByte_call_acks(0),
          dataR => accessMemoryByte_call_data(144 downto 0),
          tagR => accessMemoryByte_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryByte_return_acks(0), -- cross-over
          ackL => accessMemoryByte_return_reqs(0), -- cross-over
          dataL => accessMemoryByte_return_data(7 downto 0),
          tagL => accessMemoryByte_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity setGlobalSignals is -- 
  generic (tag_length : integer); 
  port ( -- 
    NIC_INTR_ENABLE : in std_logic_vector(0 downto 0);
    NIC_INTR_INTERNAL : in std_logic_vector(0 downto 0);
    NIC_INTR_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_INTR_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_INTR_pipe_write_data : out  std_logic_vector(0 downto 0);
    NIC_INTR_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_INTR_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_INTR_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
    S_CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    S_CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    S_CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    S_NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    S_NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    S_NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_call_acks : in   std_logic_vector(0 downto 0);
    accessRegister_call_data : out  std_logic_vector(44 downto 0);
    accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    accessRegister_return_acks : in   std_logic_vector(0 downto 0);
    accessRegister_return_data : in   std_logic_vector(31 downto 0);
    accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setGlobalSignals;
architecture setGlobalSignals_arch of setGlobalSignals is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal setGlobalSignals_CP_3610_start: Boolean;
  signal setGlobalSignals_CP_3610_symbol: Boolean;
  -- volatile/operator module components. 
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal BITSEL_u32_u1_2010_inst_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_2002_inst_req_1 : boolean;
  signal BITSEL_u32_u1_2005_inst_req_0 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_1999_inst_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_2002_inst_ack_1 : boolean;
  signal BITSEL_u32_u1_2005_inst_ack_1 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_1999_inst_ack_0 : boolean;
  signal BITSEL_u32_u1_2010_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_2013_inst_req_1 : boolean;
  signal WPIPE_NIC_INTR_2013_inst_ack_1 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_1989_inst_req_0 : boolean;
  signal BITSEL_u32_u1_2005_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2007_inst_req_1 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_1999_inst_req_1 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_1989_inst_ack_0 : boolean;
  signal call_stmt_1988_call_req_0 : boolean;
  signal call_stmt_1998_call_req_0 : boolean;
  signal WPIPE_S_CONTROL_REGISTER_1999_inst_ack_1 : boolean;
  signal call_stmt_1988_call_ack_0 : boolean;
  signal WPIPE_NIC_INTR_2013_inst_ack_0 : boolean;
  signal WPIPE_NIC_INTR_2013_inst_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_2002_inst_ack_0 : boolean;
  signal AND_u1_u1_2016_inst_ack_0 : boolean;
  signal AND_u1_u1_2016_inst_req_0 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_1989_inst_ack_1 : boolean;
  signal call_stmt_1998_call_ack_1 : boolean;
  signal BITSEL_u32_u1_2005_inst_req_1 : boolean;
  signal call_stmt_1998_call_ack_0 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2007_inst_ack_0 : boolean;
  signal BITSEL_u32_u1_2010_inst_req_1 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2007_inst_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_2002_inst_req_0 : boolean;
  signal call_stmt_1998_call_req_1 : boolean;
  signal WPIPE_S_NUMBER_OF_SERVERS_1989_inst_req_1 : boolean;
  signal BITSEL_u32_u1_2010_inst_ack_1 : boolean;
  signal AND_u1_u1_2016_inst_ack_1 : boolean;
  signal call_stmt_1988_call_ack_1 : boolean;
  signal AND_u1_u1_2016_inst_req_1 : boolean;
  signal call_stmt_1988_call_req_1 : boolean;
  signal WPIPE_NIC_INTR_ENABLE_2007_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setGlobalSignals_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setGlobalSignals_CP_3610_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setGlobalSignals_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setGlobalSignals_CP_3610_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setGlobalSignals_CP_3610_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setGlobalSignals_CP_3610_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setGlobalSignals_CP_3610: Block -- control-path 
    signal setGlobalSignals_CP_3610_elements: BooleanArray(21 downto 0);
    -- 
  begin -- 
    setGlobalSignals_CP_3610_elements(0) <= setGlobalSignals_CP_3610_start;
    setGlobalSignals_CP_3610_symbol <= setGlobalSignals_CP_3610_elements(21);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_sample_start_
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_update_start_
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/$entry
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Sample/crr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Update/ccr
      -- CP-element group 0: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Update/$entry
      -- 
    crr_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(0), ack => call_stmt_1988_call_req_0); -- 
    ccr_3628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(0), ack => call_stmt_1988_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_sample_completed_
      -- CP-element group 1: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Sample/cra
      -- 
    cra_3624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1988_call_ack_0, ack => setGlobalSignals_CP_3610_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_update_completed_
      -- CP-element group 2: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Sample/req
      -- CP-element group 2: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_sample_start_
      -- CP-element group 2: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Update/cca
      -- CP-element group 2: 	 call_stmt_1988_to_assign_stmt_1991/call_stmt_1988_Update/$exit
      -- 
    cca_3629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1988_call_ack_1, ack => setGlobalSignals_CP_3610_elements(2)); -- 
    req_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(2), ack => WPIPE_S_NUMBER_OF_SERVERS_1989_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Sample/ack
      -- CP-element group 3: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Update/$entry
      -- CP-element group 3: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Update/req
      -- CP-element group 3: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_update_start_
      -- CP-element group 3: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_sample_completed_
      -- 
    ack_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_NUMBER_OF_SERVERS_1989_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(3)); -- 
    req_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(3), ack => WPIPE_S_NUMBER_OF_SERVERS_1989_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	14 
    -- CP-element group 4:  members (17) 
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_sample_start_
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_update_start_
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_update_start_
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/$entry
      -- CP-element group 4: 	 call_stmt_1988_to_assign_stmt_1991/$exit
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Update/$entry
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Update/$entry
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Sample/crr
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_update_start_
      -- CP-element group 4: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Update/$exit
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Update/$entry
      -- CP-element group 4: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_Update/ack
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Update/cr
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Update/cr
      -- CP-element group 4: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Update/ccr
      -- CP-element group 4: 	 call_stmt_1988_to_assign_stmt_1991/WPIPE_S_NUMBER_OF_SERVERS_1989_update_completed_
      -- 
    ack_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_NUMBER_OF_SERVERS_1989_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(4)); -- 
    crr_3654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(4), ack => call_stmt_1998_call_req_0); -- 
    ccr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(4), ack => call_stmt_1998_call_req_1); -- 
    cr_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(4), ack => BITSEL_u32_u1_2005_inst_req_1); -- 
    cr_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(4), ack => BITSEL_u32_u1_2010_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_sample_completed_
      -- CP-element group 5: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Sample/$exit
      -- CP-element group 5: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Sample/cra
      -- 
    cra_3655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1998_call_ack_0, ack => setGlobalSignals_CP_3610_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6: 	13 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Sample/rr
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Sample/rr
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Sample/req
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_update_completed_
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_sample_start_
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Update/$exit
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_sample_start_
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_sample_start_
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1998_to_assign_stmt_2011/call_stmt_1998_Update/cca
      -- 
    cca_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1998_call_ack_1, ack => setGlobalSignals_CP_3610_elements(6)); -- 
    req_3668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(6), ack => WPIPE_S_CONTROL_REGISTER_1999_inst_req_0); -- 
    rr_3682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(6), ack => BITSEL_u32_u1_2005_inst_req_0); -- 
    rr_3710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(6), ack => BITSEL_u32_u1_2010_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_update_start_
      -- CP-element group 7: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Sample/$exit
      -- CP-element group 7: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Sample/ack
      -- CP-element group 7: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Update/$entry
      -- CP-element group 7: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Update/req
      -- CP-element group 7: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_sample_completed_
      -- 
    ack_3669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_CONTROL_REGISTER_1999_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(7)); -- 
    req_3673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(7), ack => WPIPE_S_CONTROL_REGISTER_1999_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	17 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_update_completed_
      -- CP-element group 8: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Update/$exit
      -- CP-element group 8: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_S_CONTROL_REGISTER_1999_Update/ack
      -- 
    ack_3674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_S_CONTROL_REGISTER_1999_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Sample/ra
      -- CP-element group 9: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_sample_completed_
      -- CP-element group 9: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Sample/$exit
      -- 
    ra_3683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u32_u1_2005_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Update/ca
      -- CP-element group 10: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_sample_start_
      -- CP-element group 10: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_update_completed_
      -- CP-element group 10: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2005_Update/$exit
      -- CP-element group 10: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Sample/req
      -- CP-element group 10: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Sample/$entry
      -- 
    ca_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u32_u1_2005_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(10)); -- 
    req_3696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(10), ack => WPIPE_MAC_ENABLE_2002_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Update/req
      -- CP-element group 11: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_sample_completed_
      -- CP-element group 11: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_update_start_
      -- CP-element group 11: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Update/$entry
      -- CP-element group 11: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Sample/ack
      -- CP-element group 11: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Sample/$exit
      -- 
    ack_3697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_2002_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(11)); -- 
    req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(11), ack => WPIPE_MAC_ENABLE_2002_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	17 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Update/$exit
      -- CP-element group 12: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_Update/ack
      -- CP-element group 12: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_MAC_ENABLE_2002_update_completed_
      -- 
    ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_2002_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	6 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Sample/$exit
      -- CP-element group 13: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Sample/ra
      -- CP-element group 13: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_sample_completed_
      -- 
    ra_3711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u32_u1_2010_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	4 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Sample/$entry
      -- CP-element group 14: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_update_completed_
      -- CP-element group 14: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Update/$exit
      -- CP-element group 14: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Sample/req
      -- CP-element group 14: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_sample_start_
      -- CP-element group 14: 	 call_stmt_1998_to_assign_stmt_2011/BITSEL_u32_u1_2010_Update/ca
      -- 
    ca_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u32_u1_2010_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(14)); -- 
    req_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(14), ack => WPIPE_NIC_INTR_ENABLE_2007_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_update_start_
      -- CP-element group 15: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Sample/$exit
      -- CP-element group 15: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Update/req
      -- CP-element group 15: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_sample_completed_
      -- CP-element group 15: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Update/$entry
      -- CP-element group 15: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Sample/ack
      -- 
    ack_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_ENABLE_2007_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(15)); -- 
    req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(15), ack => WPIPE_NIC_INTR_ENABLE_2007_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_update_completed_
      -- CP-element group 16: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Update/$exit
      -- CP-element group 16: 	 call_stmt_1998_to_assign_stmt_2011/WPIPE_NIC_INTR_ENABLE_2007_Update/ack
      -- 
    ack_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_ENABLE_2007_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: 	12 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (8) 
      -- CP-element group 17: 	 assign_stmt_2017/$entry
      -- CP-element group 17: 	 assign_stmt_2017/AND_u1_u1_2016_update_start_
      -- CP-element group 17: 	 call_stmt_1998_to_assign_stmt_2011/$exit
      -- CP-element group 17: 	 assign_stmt_2017/AND_u1_u1_2016_Update/$entry
      -- CP-element group 17: 	 assign_stmt_2017/AND_u1_u1_2016_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_2017/AND_u1_u1_2016_Sample/rr
      -- CP-element group 17: 	 assign_stmt_2017/AND_u1_u1_2016_sample_start_
      -- CP-element group 17: 	 assign_stmt_2017/AND_u1_u1_2016_Update/cr
      -- 
    rr_3741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(17), ack => AND_u1_u1_2016_inst_req_0); -- 
    cr_3746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(17), ack => AND_u1_u1_2016_inst_req_1); -- 
    setGlobalSignals_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "setGlobalSignals_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= setGlobalSignals_CP_3610_elements(8) & setGlobalSignals_CP_3610_elements(12) & setGlobalSignals_CP_3610_elements(16);
      gj_setGlobalSignals_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => setGlobalSignals_CP_3610_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_2017/AND_u1_u1_2016_sample_completed_
      -- CP-element group 18: 	 assign_stmt_2017/AND_u1_u1_2016_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_2017/AND_u1_u1_2016_Sample/ra
      -- 
    ra_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2016_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_sample_start_
      -- CP-element group 19: 	 assign_stmt_2017/AND_u1_u1_2016_Update/$exit
      -- CP-element group 19: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Sample/req
      -- CP-element group 19: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Sample/$entry
      -- CP-element group 19: 	 assign_stmt_2017/AND_u1_u1_2016_update_completed_
      -- CP-element group 19: 	 assign_stmt_2017/AND_u1_u1_2016_Update/ca
      -- 
    ca_3747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_2016_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(19)); -- 
    req_3755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(19), ack => WPIPE_NIC_INTR_2013_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_update_start_
      -- CP-element group 20: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Update/req
      -- CP-element group 20: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Update/$entry
      -- CP-element group 20: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Sample/ack
      -- CP-element group 20: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_sample_completed_
      -- 
    ack_3756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_2013_inst_ack_0, ack => setGlobalSignals_CP_3610_elements(20)); -- 
    req_3760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setGlobalSignals_CP_3610_elements(20), ack => WPIPE_NIC_INTR_2013_inst_req_1); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 $exit
      -- CP-element group 21: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Update/$exit
      -- CP-element group 21: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_Update/ack
      -- CP-element group 21: 	 assign_stmt_2017/WPIPE_NIC_INTR_2013_update_completed_
      -- CP-element group 21: 	 assign_stmt_2017/$exit
      -- 
    ack_3761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_INTR_2013_inst_ack_1, ack => setGlobalSignals_CP_3610_elements(21)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_2016_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2005_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2010_wire : std_logic_vector(0 downto 0);
    signal RPIPE_NIC_INTR_ENABLE_2014_wire : std_logic_vector(0 downto 0);
    signal RPIPE_NIC_INTR_INTERNAL_2015_wire : std_logic_vector(0 downto 0);
    signal R_READMEM_1983_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_1993_wire_constant : std_logic_vector(0 downto 0);
    signal ctrl_reg_1998 : std_logic_vector(31 downto 0);
    signal konst_1984_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1985_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1986_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1994_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1995_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1996_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2004_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2009_wire_constant : std_logic_vector(31 downto 0);
    signal n_servers_1988 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_READMEM_1983_wire_constant <= "1";
    R_READMEM_1993_wire_constant <= "1";
    konst_1984_wire_constant <= "1111";
    konst_1985_wire_constant <= "00000001";
    konst_1986_wire_constant <= "00000000000000000000000000000000";
    konst_1994_wire_constant <= "1111";
    konst_1995_wire_constant <= "00000000";
    konst_1996_wire_constant <= "00000000000000000000000000000000";
    konst_2004_wire_constant <= "00000000000000000000000000000001";
    konst_2009_wire_constant <= "00000000000000000000000000000010";
    -- shared split operator group (0) : AND_u1_u1_2016_inst 
    ApIntAnd_group_0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_NIC_INTR_ENABLE_2014_wire & RPIPE_NIC_INTR_INTERNAL_2015_wire;
      AND_u1_u1_2016_wire <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_2016_inst_req_0;
      AND_u1_u1_2016_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_2016_inst_req_1;
      AND_u1_u1_2016_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : BITSEL_u32_u1_2005_inst 
    ApBitsel_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ctrl_reg_1998;
      BITSEL_u32_u1_2005_wire <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u32_u1_2005_inst_req_0;
      BITSEL_u32_u1_2005_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u32_u1_2005_inst_req_1;
      BITSEL_u32_u1_2005_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_1_gI: SplitGuardInterface generic map(name => "ApBitsel_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : BITSEL_u32_u1_2010_inst 
    ApBitsel_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ctrl_reg_1998;
      BITSEL_u32_u1_2010_wire <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u32_u1_2010_inst_req_0;
      BITSEL_u32_u1_2010_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u32_u1_2010_inst_req_1;
      BITSEL_u32_u1_2010_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_2_gI: SplitGuardInterface generic map(name => "ApBitsel_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- read from input-signal NIC_INTR_ENABLE
    RPIPE_NIC_INTR_ENABLE_2014_wire <= NIC_INTR_ENABLE;
    -- read from input-signal NIC_INTR_INTERNAL
    RPIPE_NIC_INTR_INTERNAL_2015_wire <= NIC_INTR_INTERNAL;
    -- shared outport operator group (0) : WPIPE_MAC_ENABLE_2002_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_MAC_ENABLE_2002_inst_req_0;
      WPIPE_MAC_ENABLE_2002_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_MAC_ENABLE_2002_inst_req_1;
      WPIPE_MAC_ENABLE_2002_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= BITSEL_u32_u1_2005_wire;
      MAC_ENABLE_write_0_gI: SplitGuardInterface generic map(name => "MAC_ENABLE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      MAC_ENABLE_write_0: OutputPortRevised -- 
        generic map ( name => "MAC_ENABLE", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => MAC_ENABLE_pipe_write_req(0),
          oack => MAC_ENABLE_pipe_write_ack(0),
          odata => MAC_ENABLE_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_NIC_INTR_2013_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_INTR_2013_inst_req_0;
      WPIPE_NIC_INTR_2013_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_INTR_2013_inst_req_1;
      WPIPE_NIC_INTR_2013_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= AND_u1_u1_2016_wire;
      NIC_INTR_write_1_gI: SplitGuardInterface generic map(name => "NIC_INTR_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_INTR_write_1: OutputPortRevised -- 
        generic map ( name => "NIC_INTR", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_INTR_pipe_write_req(0),
          oack => NIC_INTR_pipe_write_ack(0),
          odata => NIC_INTR_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_NIC_INTR_ENABLE_2007_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_INTR_ENABLE_2007_inst_req_0;
      WPIPE_NIC_INTR_ENABLE_2007_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_INTR_ENABLE_2007_inst_req_1;
      WPIPE_NIC_INTR_ENABLE_2007_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= BITSEL_u32_u1_2010_wire;
      NIC_INTR_ENABLE_write_2_gI: SplitGuardInterface generic map(name => "NIC_INTR_ENABLE_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_INTR_ENABLE_write_2: OutputPortRevised -- 
        generic map ( name => "NIC_INTR_ENABLE", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_INTR_ENABLE_pipe_write_req(0),
          oack => NIC_INTR_ENABLE_pipe_write_ack(0),
          odata => NIC_INTR_ENABLE_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_S_CONTROL_REGISTER_1999_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_S_CONTROL_REGISTER_1999_inst_req_0;
      WPIPE_S_CONTROL_REGISTER_1999_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_S_CONTROL_REGISTER_1999_inst_req_1;
      WPIPE_S_CONTROL_REGISTER_1999_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= ctrl_reg_1998;
      S_CONTROL_REGISTER_write_3_gI: SplitGuardInterface generic map(name => "S_CONTROL_REGISTER_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      S_CONTROL_REGISTER_write_3: OutputPortRevised -- 
        generic map ( name => "S_CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => S_CONTROL_REGISTER_pipe_write_req(0),
          oack => S_CONTROL_REGISTER_pipe_write_ack(0),
          odata => S_CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_S_NUMBER_OF_SERVERS_1989_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_S_NUMBER_OF_SERVERS_1989_inst_req_0;
      WPIPE_S_NUMBER_OF_SERVERS_1989_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_S_NUMBER_OF_SERVERS_1989_inst_req_1;
      WPIPE_S_NUMBER_OF_SERVERS_1989_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= n_servers_1988;
      S_NUMBER_OF_SERVERS_write_4_gI: SplitGuardInterface generic map(name => "S_NUMBER_OF_SERVERS_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      S_NUMBER_OF_SERVERS_write_4: OutputPortRevised -- 
        generic map ( name => "S_NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => S_NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => S_NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => S_NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1988_call call_stmt_1998_call 
    accessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(89 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1988_call_req_0;
      reqL_unguarded(0) <= call_stmt_1998_call_req_0;
      call_stmt_1988_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1998_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1988_call_req_1;
      reqR_unguarded(0) <= call_stmt_1998_call_req_1;
      call_stmt_1988_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1998_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "accessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_READMEM_1983_wire_constant & konst_1984_wire_constant & konst_1985_wire_constant & konst_1986_wire_constant & R_READMEM_1993_wire_constant & konst_1994_wire_constant & konst_1995_wire_constant & konst_1996_wire_constant;
      n_servers_1988 <= data_out(63 downto 32);
      ctrl_reg_1998 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 90,
        owidth => 45,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessRegister_call_reqs(0),
          ackR => accessRegister_call_acks(0),
          dataR => accessRegister_call_data(44 downto 0),
          tagR => accessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessRegister_return_acks(0), -- cross-over
          ackL => accessRegister_return_reqs(0), -- cross-over
          dataL => accessRegister_return_data(31 downto 0),
          tagL => accessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setGlobalSignals_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    buf_base_address : in  std_logic_vector(63 downto 0);
    write_index : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(63 downto 0);
    accessQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueElement_call_data : out  std_logic_vector(168 downto 0);
    accessQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueElement_return_data : in   std_logic_vector(63 downto 0);
    accessQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 168)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal buf_base_address_buffer :  std_logic_vector(63 downto 0);
  signal buf_base_address_update_enable: Boolean;
  signal write_index_buffer :  std_logic_vector(31 downto 0);
  signal write_index_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(63 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_2409_start: Boolean;
  signal setQueueElement_CP_2409_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      index : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1572_call_req_1 : boolean;
  signal call_stmt_1572_call_ack_1 : boolean;
  signal call_stmt_1572_call_ack_0 : boolean;
  signal call_stmt_1572_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 168) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= buf_base_address;
  buf_base_address_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(103 downto 72) <= write_index;
  write_index_buffer <= in_buffer_data_out(103 downto 72);
  in_buffer_data_in(167 downto 104) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(167 downto 104);
  in_buffer_data_in(tag_length + 167 downto 168) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 167 downto 168);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_2409_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_2409_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_2409_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_2409_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_2409: Block -- control-path 
    signal setQueueElement_CP_2409_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_2409_elements(0) <= setQueueElement_CP_2409_start;
    setQueueElement_CP_2409_symbol <= setQueueElement_CP_2409_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_1572/call_stmt_1572_Update/$entry
      -- CP-element group 0: 	 call_stmt_1572/call_stmt_1572_Update/ccr
      -- CP-element group 0: 	 call_stmt_1572/call_stmt_1572_sample_start_
      -- CP-element group 0: 	 call_stmt_1572/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1572/call_stmt_1572_Sample/crr
      -- CP-element group 0: 	 call_stmt_1572/call_stmt_1572_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1572/call_stmt_1572_update_start_
      -- 
    crr_2422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_2409_elements(0), ack => call_stmt_1572_call_req_0); -- 
    ccr_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_2409_elements(0), ack => call_stmt_1572_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1572/call_stmt_1572_Sample/cra
      -- CP-element group 1: 	 call_stmt_1572/call_stmt_1572_sample_completed_
      -- CP-element group 1: 	 call_stmt_1572/call_stmt_1572_Sample/$exit
      -- 
    cra_2423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1572_call_ack_0, ack => setQueueElement_CP_2409_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_1572/$exit
      -- CP-element group 2: 	 call_stmt_1572/call_stmt_1572_Update/$exit
      -- CP-element group 2: 	 call_stmt_1572/call_stmt_1572_Update/cca
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1572/call_stmt_1572_update_completed_
      -- 
    cca_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1572_call_ack_1, ack => setQueueElement_CP_2409_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_WRITEMEM_1567_wire_constant : std_logic_vector(0 downto 0);
    signal q_r_data_1572 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    R_WRITEMEM_1567_wire_constant <= "0";
    -- shared call operator group (0) : call_stmt_1572_call 
    accessQueueElement_call_group_0: Block -- 
      signal data_in: std_logic_vector(168 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1572_call_req_0;
      call_stmt_1572_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1572_call_req_1;
      call_stmt_1572_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueElement_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueElement_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_WRITEMEM_1567_wire_constant & buf_base_address_buffer & write_index_buffer & q_w_data_buffer;
      q_r_data_1572 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 169,
        owidth => 169,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueElement_call_reqs(0),
          ackR => accessQueueElement_call_acks(0),
          dataR => accessQueueElement_call_data(168 downto 0),
          tagR => accessQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueElement_return_acks(0), -- cross-over
          ackL => accessQueueElement_return_reqs(0), -- cross-over
          dataL => accessQueueElement_return_data(63 downto 0),
          tagL => accessQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    q_base_address : in  std_logic_vector(63 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
    accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
    accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
    accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
    accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
    accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 136)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(63 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_1557_start: Boolean;
  signal setQueuePointers_CP_1557_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueReadIndex is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessQueueWriteIndex is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1144_call_ack_1 : boolean;
  signal call_stmt_1144_call_ack_0 : boolean;
  signal call_stmt_1144_call_req_1 : boolean;
  signal call_stmt_1144_call_req_0 : boolean;
  signal call_stmt_1150_call_req_0 : boolean;
  signal call_stmt_1150_call_ack_1 : boolean;
  signal call_stmt_1150_call_req_1 : boolean;
  signal call_stmt_1150_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 136) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(103 downto 72) <= wp;
  wp_buffer <= in_buffer_data_out(103 downto 72);
  in_buffer_data_in(135 downto 104) <= rp;
  rp_buffer <= in_buffer_data_out(135 downto 104);
  in_buffer_data_in(tag_length + 135 downto 136) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 135 downto 136);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_1557_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_1557_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_1557_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_1557_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_1557: Block -- control-path 
    signal setQueuePointers_CP_1557_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_1557_elements(0) <= setQueuePointers_CP_1557_start;
    setQueuePointers_CP_1557_symbol <= setQueuePointers_CP_1557_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_update_start_
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Update/$entry
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/$entry
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_sample_start_
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Sample/crr
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Update/ccr
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_update_start_
      -- CP-element group 0: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Update/$entry
      -- 
    crr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1557_elements(0), ack => call_stmt_1144_call_req_0); -- 
    ccr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1557_elements(0), ack => call_stmt_1144_call_req_1); -- 
    ccr_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1557_elements(0), ack => call_stmt_1150_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Sample/cra
      -- CP-element group 1: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_sample_completed_
      -- 
    cra_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1144_call_ack_0, ack => setQueuePointers_CP_1557_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Update/cca
      -- CP-element group 2: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_Update/$exit
      -- CP-element group 2: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Sample/crr
      -- CP-element group 2: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_sample_start_
      -- CP-element group 2: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1144_update_completed_
      -- 
    cca_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1144_call_ack_1, ack => setQueuePointers_CP_1557_elements(2)); -- 
    crr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1557_elements(2), ack => call_stmt_1150_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_sample_completed_
      -- CP-element group 3: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Sample/cra
      -- 
    cra_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1150_call_ack_0, ack => setQueuePointers_CP_1557_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_update_completed_
      -- CP-element group 4: 	 call_stmt_1144_to_call_stmt_1150/$exit
      -- CP-element group 4: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Update/cca
      -- CP-element group 4: 	 call_stmt_1144_to_call_stmt_1150/call_stmt_1150_Update/$exit
      -- 
    cca_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1150_call_ack_1, ack => setQueuePointers_CP_1557_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_WRITEMEM_1140_wire_constant : std_logic_vector(0 downto 0);
    signal R_WRITEMEM_1146_wire_constant : std_logic_vector(0 downto 0);
    signal ign_rp_1144 : std_logic_vector(31 downto 0);
    signal ign_wp_1150 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_WRITEMEM_1140_wire_constant <= "0";
    R_WRITEMEM_1146_wire_constant <= "0";
    -- shared call operator group (0) : call_stmt_1144_call 
    accessQueueReadIndex_call_group_0: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1144_call_req_0;
      call_stmt_1144_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1144_call_req_1;
      call_stmt_1144_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueReadIndex_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueReadIndex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_WRITEMEM_1140_wire_constant & q_base_address_buffer & rp_buffer;
      ign_rp_1144 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueReadIndex_call_reqs(0),
          ackR => accessQueueReadIndex_call_acks(0),
          dataR => accessQueueReadIndex_call_data(104 downto 0),
          tagR => accessQueueReadIndex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueReadIndex_return_acks(0), -- cross-over
          ackL => accessQueueReadIndex_return_reqs(0), -- cross-over
          dataL => accessQueueReadIndex_return_data(31 downto 0),
          tagL => accessQueueReadIndex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1150_call 
    accessQueueWriteIndex_call_group_1: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1150_call_req_0;
      call_stmt_1150_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1150_call_req_1;
      call_stmt_1150_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueWriteIndex_call_group_1_gI: SplitGuardInterface generic map(name => "accessQueueWriteIndex_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_WRITEMEM_1146_wire_constant & q_base_address_buffer & wp_buffer;
      ign_wp_1150 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueWriteIndex_call_reqs(0),
          ackR => accessQueueWriteIndex_call_acks(0),
          dataR => accessQueueWriteIndex_call_data(104 downto 0),
          tagR => accessQueueWriteIndex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueWriteIndex_return_acks(0), -- cross-over
          ackL => accessQueueWriteIndex_return_reqs(0), -- cross-over
          dataL => accessQueueWriteIndex_return_data(31 downto 0),
          tagL => accessQueueWriteIndex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity setTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    q_base_address : in  std_logic_vector(63 downto 0);
    updated_total_msgs : in  std_logic_vector(31 downto 0);
    accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
    accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
    accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
    accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setTotalMessages;
architecture setTotalMessages_arch of setTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(63 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal updated_total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal updated_total_msgs_update_enable: Boolean;
  -- output port buffer signals
  signal setTotalMessages_CP_1591_start: Boolean;
  signal setTotalMessages_CP_1591_symbol: Boolean;
  -- volatile/operator module components. 
  component accessQueueTotalMsgs is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1161_call_ack_1 : boolean;
  signal call_stmt_1161_call_req_1 : boolean;
  signal call_stmt_1161_call_ack_0 : boolean;
  signal call_stmt_1161_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(103 downto 72) <= updated_total_msgs;
  updated_total_msgs_buffer <= in_buffer_data_out(103 downto 72);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setTotalMessages_CP_1591_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setTotalMessages_CP_1591_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setTotalMessages_CP_1591_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setTotalMessages_CP_1591_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setTotalMessages_CP_1591: Block -- control-path 
    signal setTotalMessages_CP_1591_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setTotalMessages_CP_1591_elements(0) <= setTotalMessages_CP_1591_start;
    setTotalMessages_CP_1591_symbol <= setTotalMessages_CP_1591_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1161/call_stmt_1161_sample_start_
      -- CP-element group 0: 	 call_stmt_1161/$entry
      -- CP-element group 0: 	 call_stmt_1161/call_stmt_1161_Update/ccr
      -- CP-element group 0: 	 call_stmt_1161/call_stmt_1161_Update/$entry
      -- CP-element group 0: 	 call_stmt_1161/call_stmt_1161_Sample/crr
      -- CP-element group 0: 	 call_stmt_1161/call_stmt_1161_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1161/call_stmt_1161_update_start_
      -- 
    ccr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setTotalMessages_CP_1591_elements(0), ack => call_stmt_1161_call_req_1); -- 
    crr_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setTotalMessages_CP_1591_elements(0), ack => call_stmt_1161_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1161/call_stmt_1161_sample_completed_
      -- CP-element group 1: 	 call_stmt_1161/call_stmt_1161_Sample/cra
      -- CP-element group 1: 	 call_stmt_1161/call_stmt_1161_Sample/$exit
      -- 
    cra_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1161_call_ack_0, ack => setTotalMessages_CP_1591_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1161/call_stmt_1161_Update/cca
      -- CP-element group 2: 	 call_stmt_1161/$exit
      -- CP-element group 2: 	 call_stmt_1161/call_stmt_1161_Update/$exit
      -- CP-element group 2: 	 call_stmt_1161/call_stmt_1161_update_completed_
      -- 
    cca_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1161_call_ack_1, ack => setTotalMessages_CP_1591_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_WRITEMEM_1157_wire_constant : std_logic_vector(0 downto 0);
    signal ignore_1161 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_WRITEMEM_1157_wire_constant <= "0";
    -- shared call operator group (0) : call_stmt_1161_call 
    accessQueueTotalMsgs_call_group_0: Block -- 
      signal data_in: std_logic_vector(104 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1161_call_req_0;
      call_stmt_1161_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1161_call_req_1;
      call_stmt_1161_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessQueueTotalMsgs_call_group_0_gI: SplitGuardInterface generic map(name => "accessQueueTotalMsgs_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_WRITEMEM_1157_wire_constant & q_base_address_buffer & updated_total_msgs_buffer;
      ignore_1161 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 105,
        owidth => 105,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessQueueTotalMsgs_call_reqs(0),
          ackR => accessQueueTotalMsgs_call_acks(0),
          dataR => accessQueueTotalMsgs_call_data(104 downto 0),
          tagR => accessQueueTotalMsgs_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessQueueTotalMsgs_return_acks(0), -- cross-over
          ackL => accessQueueTotalMsgs_return_reqs(0), -- cross-over
          dataL => accessQueueTotalMsgs_return_data(31 downto 0),
          tagL => accessQueueTotalMsgs_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(7 downto 0);
    S_CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    S_NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(15 downto 0);
    TX_ACTIVITY_LOGGER_pipe_write_req : out  std_logic_vector(0 downto 0);
    TX_ACTIVITY_LOGGER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    TX_ACTIVITY_LOGGER_pipe_write_data : out  std_logic_vector(7 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(15 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(64 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    incrementNumberOfPacketsTransmitted_call_reqs : out  std_logic_vector(0 downto 0);
    incrementNumberOfPacketsTransmitted_call_acks : in   std_logic_vector(0 downto 0);
    incrementNumberOfPacketsTransmitted_call_tag  :  out  std_logic_vector(0 downto 0);
    incrementNumberOfPacketsTransmitted_return_reqs : out  std_logic_vector(0 downto 0);
    incrementNumberOfPacketsTransmitted_return_acks : in   std_logic_vector(0 downto 0);
    incrementNumberOfPacketsTransmitted_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(71 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_4738_start: Boolean;
  signal transmitEngineDaemon_CP_4738_symbol: Boolean;
  -- volatile/operator module components. 
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_w_data : in  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(167 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      server_index : in  std_logic_vector(7 downto 0);
      pkt_pointer : out  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(17 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(64 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component incrementNumberOfPacketsTransmitted is -- 
    generic (tag_length : integer); 
    port ( -- 
      incrementRegister_call_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_call_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_call_data : out  std_logic_vector(7 downto 0);
      incrementRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementRegister_return_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_return_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_return_data : in   std_logic_vector(31 downto 0);
      incrementRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      packet_pointer : in  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(1 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(401 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(1 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(127 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_ack_1 : boolean;
  signal if_stmt_2511_branch_req_0 : boolean;
  signal if_stmt_2511_branch_ack_1 : boolean;
  signal if_stmt_2511_branch_ack_0 : boolean;
  signal do_while_stmt_2522_branch_req_0 : boolean;
  signal AND_u8_u8_2533_inst_req_0 : boolean;
  signal AND_u8_u8_2533_inst_ack_0 : boolean;
  signal AND_u8_u8_2533_inst_req_1 : boolean;
  signal AND_u8_u8_2533_inst_ack_1 : boolean;
  signal phi_stmt_2534_req_0 : boolean;
  signal phi_stmt_2534_req_1 : boolean;
  signal phi_stmt_2534_ack_0 : boolean;
  signal call_stmt_2547_call_req_0 : boolean;
  signal call_stmt_2547_call_ack_0 : boolean;
  signal call_stmt_2547_call_req_1 : boolean;
  signal call_stmt_2547_call_ack_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2549_inst_req_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2549_inst_ack_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2549_inst_req_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2549_inst_ack_1 : boolean;
  signal call_stmt_2556_call_req_0 : boolean;
  signal call_stmt_2556_call_ack_0 : boolean;
  signal call_stmt_2556_call_req_1 : boolean;
  signal call_stmt_2556_call_ack_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2558_inst_req_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2558_inst_ack_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2558_inst_req_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2558_inst_ack_1 : boolean;
  signal NOT_u1_u1_2563_inst_req_0 : boolean;
  signal NOT_u1_u1_2563_inst_ack_0 : boolean;
  signal NOT_u1_u1_2563_inst_req_1 : boolean;
  signal NOT_u1_u1_2563_inst_ack_1 : boolean;
  signal W_pkt_pointer_2477_delayed_4_0_2573_inst_req_0 : boolean;
  signal W_pkt_pointer_2477_delayed_4_0_2573_inst_ack_0 : boolean;
  signal W_pkt_pointer_2477_delayed_4_0_2573_inst_req_1 : boolean;
  signal W_pkt_pointer_2477_delayed_4_0_2573_inst_ack_1 : boolean;
  signal call_stmt_2582_call_req_0 : boolean;
  signal call_stmt_2582_call_ack_0 : boolean;
  signal call_stmt_2582_call_req_1 : boolean;
  signal call_stmt_2582_call_ack_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2584_inst_req_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2584_inst_ack_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2584_inst_req_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2584_inst_ack_1 : boolean;
  signal call_stmt_2590_call_req_0 : boolean;
  signal call_stmt_2590_call_ack_0 : boolean;
  signal call_stmt_2590_call_req_1 : boolean;
  signal call_stmt_2590_call_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_ack_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2595_inst_req_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2595_inst_ack_0 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2595_inst_req_1 : boolean;
  signal WPIPE_TX_ACTIVITY_LOGGER_2595_inst_ack_1 : boolean;
  signal do_while_stmt_2522_branch_ack_0 : boolean;
  signal do_while_stmt_2522_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_4738_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_4738_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_4738_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_4738_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_4738: Block -- control-path 
    signal transmitEngineDaemon_CP_4738_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_4738_elements(0) <= transmitEngineDaemon_CP_4738_start;
    transmitEngineDaemon_CP_4738_symbol <= transmitEngineDaemon_CP_4738_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_2508/$entry
      -- CP-element group 0: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_sample_start_
      -- CP-element group 0: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Sample/req
      -- 
    req_4751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_sample_completed_
      -- CP-element group 1: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_update_start_
      -- CP-element group 1: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Sample/ack
      -- CP-element group 1: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Update/$entry
      -- CP-element group 1: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Update/req
      -- 
    ack_4752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(1)); -- 
    req_4756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	89 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_2508/$exit
      -- CP-element group 2: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_update_completed_
      -- CP-element group 2: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Update/$exit
      -- CP-element group 2: 	 assign_stmt_2508/WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_2509/$entry
      -- CP-element group 2: 	 branch_block_stmt_2509/branch_block_stmt_2509__entry__
      -- CP-element group 2: 	 branch_block_stmt_2509/merge_stmt_2510__entry__
      -- CP-element group 2: 	 branch_block_stmt_2509/merge_stmt_2510_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_2509/merge_stmt_2510__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_2509/merge_stmt_2510__entry___PhiReq/$exit
      -- 
    ack_4757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_2509/$exit
      -- CP-element group 3: 	 branch_block_stmt_2509/branch_block_stmt_2509__exit__
      -- 
    transmitEngineDaemon_CP_4738_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	88 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	89 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_2509/do_while_stmt_2522__exit__
      -- CP-element group 4: 	 branch_block_stmt_2509/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_2509/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_2509/disable_loopback_PhiReq/$exit
      -- 
    transmitEngineDaemon_CP_4738_elements(4) <= transmitEngineDaemon_CP_4738_elements(88);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	89 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	89 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2509/if_stmt_2511_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_2509/if_stmt_2511_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_2509/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_2509/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_2509/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_4832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2511_branch_ack_1, ack => transmitEngineDaemon_CP_4738_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	89 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (8) 
      -- CP-element group 6: 	 branch_block_stmt_2509/if_stmt_2511__exit__
      -- CP-element group 6: 	 branch_block_stmt_2509/assign_stmt_2520__entry__
      -- CP-element group 6: 	 branch_block_stmt_2509/assign_stmt_2520__exit__
      -- CP-element group 6: 	 branch_block_stmt_2509/do_while_stmt_2522__entry__
      -- CP-element group 6: 	 branch_block_stmt_2509/if_stmt_2511_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_2509/if_stmt_2511_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_2509/assign_stmt_2520/$entry
      -- CP-element group 6: 	 branch_block_stmt_2509/assign_stmt_2520/$exit
      -- 
    else_choice_transition_4836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2511_branch_ack_0, ack => transmitEngineDaemon_CP_4738_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_2509/do_while_stmt_2522/$entry
      -- CP-element group 7: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522__entry__
      -- 
    transmitEngineDaemon_CP_4738_elements(7) <= transmitEngineDaemon_CP_4738_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	88 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522__exit__
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_back
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	86 
    -- CP-element group 10: 	87 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2509/do_while_stmt_2522/condition_done
      -- CP-element group 10: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_taken/$entry
      -- 
    transmitEngineDaemon_CP_4738_elements(10) <= transmitEngineDaemon_CP_4738_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	85 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_body_done
      -- 
    transmitEngineDaemon_CP_4738_elements(11) <= transmitEngineDaemon_CP_4738_elements(85);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	30 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/back_edge_to_loop_body
      -- 
    transmitEngineDaemon_CP_4738_elements(12) <= transmitEngineDaemon_CP_4738_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	32 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/first_time_through_loop_body
      -- 
    transmitEngineDaemon_CP_4738_elements(13) <= transmitEngineDaemon_CP_4738_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	82 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	27 
    -- CP-element group 14: 	26 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2524_sample_start_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	82 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/condition_evaluated
      -- 
    condition_evaluated_4855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(15), ack => do_while_stmt_2522_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(20) & transmitEngineDaemon_CP_4738_elements(82);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	26 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_sample_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(14) & transmitEngineDaemon_CP_4738_elements(26) & transmitEngineDaemon_CP_4738_elements(20);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	28 
    -- CP-element group 17: 	24 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	85 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	26 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2524_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_sample_completed_
      -- 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(28) & transmitEngineDaemon_CP_4738_elements(24);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	85 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(18) is a control-delay.
    cp_element_18_delay: control_delay_element  generic map(name => " 18_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_4738_elements(17), ack => transmitEngineDaemon_CP_4738_elements(18), clk => clk, reset =>reset);
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	27 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/aggregated_phi_update_req
      -- CP-element group 19: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_update_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(21) & transmitEngineDaemon_CP_4738_elements(27);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	29 
    -- CP-element group 20: 	25 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/aggregated_phi_update_ack
      -- 
    transmitEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(29) & transmitEngineDaemon_CP_4738_elements(25);
      gj_transmitEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	77 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2524_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(14) & transmitEngineDaemon_CP_4738_elements(45) & transmitEngineDaemon_CP_4738_elements(77);
      gj_transmitEngineDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Sample/rr
      -- 
    rr_4873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(22), ack => AND_u8_u8_2533_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(16) & transmitEngineDaemon_CP_4738_elements(24);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_update_start_
      -- CP-element group 23: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Update/cr
      -- 
    cr_4878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(23), ack => AND_u8_u8_2533_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(19) & transmitEngineDaemon_CP_4738_elements(25);
      gj_transmitEngineDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Sample/ra
      -- 
    ra_4874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u8_u8_2533_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	43 
    -- CP-element group 25: 	76 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2524_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/AND_u8_u8_2533_Update/ca
      -- 
    ca_4879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u8_u8_2533_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	16 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_sample_start_
      -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(14) & transmitEngineDaemon_CP_4738_elements(17);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	19 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(14) & transmitEngineDaemon_CP_4738_elements(29);
      gj_transmitEngineDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	17 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_sample_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	20 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_update_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	12 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_loopback_trigger
      -- 
    transmitEngineDaemon_CP_4738_elements(30) <= transmitEngineDaemon_CP_4738_elements(12);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_loopback_sample_req
      -- CP-element group 31: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_loopback_sample_req_ps
      -- 
    phi_stmt_2534_loopback_sample_req_4889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2534_loopback_sample_req_4889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(31), ack => phi_stmt_2534_req_0); -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	13 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_entry_trigger
      -- 
    transmitEngineDaemon_CP_4738_elements(32) <= transmitEngineDaemon_CP_4738_elements(13);
    -- CP-element group 33:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_entry_sample_req
      -- CP-element group 33: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_entry_sample_req_ps
      -- 
    phi_stmt_2534_entry_sample_req_4892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2534_entry_sample_req_4892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(33), ack => phi_stmt_2534_req_1); -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_phi_mux_ack
      -- CP-element group 34: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/phi_stmt_2534_phi_mux_ack_ps
      -- 
    phi_stmt_2534_phi_mux_ack_4895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2534_ack_0, ack => transmitEngineDaemon_CP_4738_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_sample_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_update_start_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_update_completed__ps
      -- 
    transmitEngineDaemon_CP_4738_elements(37) <= transmitEngineDaemon_CP_4738_elements(38);
    -- CP-element group 38:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	37 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2537_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_4738_elements(36), ack => transmitEngineDaemon_CP_4738_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_sample_start__ps
      -- CP-element group 39: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_sample_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_update_start__ps
      -- CP-element group 40: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_update_start_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_update_completed__ps
      -- 
    transmitEngineDaemon_CP_4738_elements(41) <= transmitEngineDaemon_CP_4738_elements(42);
    -- CP-element group 42:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	41 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/type_cast_2539_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(42) is a control-delay.
    cp_element_42_delay: control_delay_element  generic map(name => " 42_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_4738_elements(40), ack => transmitEngineDaemon_CP_4738_elements(42), clk => clk, reset =>reset);
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	25 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	67 
    -- CP-element group 43: 	75 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Sample/crr
      -- 
    crr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(43), ack => call_stmt_2547_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(25) & transmitEngineDaemon_CP_4738_elements(67) & transmitEngineDaemon_CP_4738_elements(75);
      gj_transmitEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	62 
    -- CP-element group 44: 	51 
    -- CP-element group 44: 	58 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_update_start_
      -- CP-element group 44: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Update/ccr
      -- 
    ccr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(44), ack => call_stmt_2547_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(62) & transmitEngineDaemon_CP_4738_elements(51) & transmitEngineDaemon_CP_4738_elements(58);
      gj_transmitEngineDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	21 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Sample/cra
      -- 
    cra_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2547_call_ack_0, ack => transmitEngineDaemon_CP_4738_elements(45)); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	83 
    -- CP-element group 46: 	51 
    -- CP-element group 46: 	60 
    -- CP-element group 46:  members (7) 
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_Update/cca
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/barrier_stmt_2548_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Sample/crr
      -- 
    cca_4927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2547_call_ack_1, ack => transmitEngineDaemon_CP_4738_elements(46)); -- 
    crr_4950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(46), ack => call_stmt_2556_call_req_0); -- 
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	81 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Sample/req
      -- 
    req_4936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(47), ack => WPIPE_TX_ACTIVITY_LOGGER_2549_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(46) & transmitEngineDaemon_CP_4738_elements(81);
      gj_transmitEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_update_start_
      -- CP-element group 48: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Update/req
      -- 
    ack_4937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2549_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(48)); -- 
    req_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(48), ack => WPIPE_TX_ACTIVITY_LOGGER_2549_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	53 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2549_Update/ack
      -- 
    ack_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2549_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	66 
    -- CP-element group 50: 	74 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_update_start_
      -- CP-element group 50: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Update/ccr
      -- 
    ccr_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(50), ack => call_stmt_2556_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(66) & transmitEngineDaemon_CP_4738_elements(74);
      gj_transmitEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	46 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	44 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Sample/cra
      -- 
    cra_4951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2556_call_ack_0, ack => transmitEngineDaemon_CP_4738_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	64 
    -- CP-element group 52: 	72 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2556_Update/cca
      -- 
    cca_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2556_call_ack_1, ack => transmitEngineDaemon_CP_4738_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	49 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	58 
    -- CP-element group 53: 	60 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/barrier_stmt_2557_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Sample/rr
      -- 
    rr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(53), ack => NOT_u1_u1_2563_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(49) & transmitEngineDaemon_CP_4738_elements(52);
      gj_transmitEngineDaemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Sample/req
      -- 
    req_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(54), ack => WPIPE_TX_ACTIVITY_LOGGER_2558_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(53) & transmitEngineDaemon_CP_4738_elements(56);
      gj_transmitEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Update/req
      -- 
    ack_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2558_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(55)); -- 
    req_4970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(55), ack => WPIPE_TX_ACTIVITY_LOGGER_2558_inst_req_1); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	68 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2558_Update/ack
      -- 
    ack_4971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2558_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	66 
    -- CP-element group 57: 	74 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Update/cr
      -- 
    cr_4984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(57), ack => NOT_u1_u1_2563_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(66) & transmitEngineDaemon_CP_4738_elements(74);
      gj_transmitEngineDaemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	53 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	44 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Sample/ra
      -- 
    ra_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_2563_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59: 	64 
    -- CP-element group 59: 	72 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/NOT_u1_u1_2563_Update/ca
      -- 
    ca_4985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_2563_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	46 
    -- CP-element group 60: 	53 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Sample/req
      -- 
    req_4993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(60), ack => W_pkt_pointer_2477_delayed_4_0_2573_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(46) & transmitEngineDaemon_CP_4738_elements(53);
      gj_transmitEngineDaemon_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	66 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_update_start_
      -- CP-element group 61: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Update/req
      -- 
    req_4998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(61), ack => W_pkt_pointer_2477_delayed_4_0_2573_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_4738_elements(66);
      gj_transmitEngineDaemon_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	44 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Sample/ack
      -- 
    ack_4994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_2477_delayed_4_0_2573_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/assign_stmt_2575_Update/ack
      -- 
    ack_4999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_2477_delayed_4_0_2573_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: 	83 
    -- CP-element group 64: 	52 
    -- CP-element group 64: 	59 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Sample/crr
      -- 
    crr_5007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(64), ack => call_stmt_2582_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(63) & transmitEngineDaemon_CP_4738_elements(83) & transmitEngineDaemon_CP_4738_elements(52) & transmitEngineDaemon_CP_4738_elements(59);
      gj_transmitEngineDaemon_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Update/ccr
      -- 
    ccr_5012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(65), ack => call_stmt_2582_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_4738_elements(67);
      gj_transmitEngineDaemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	61 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Sample/cra
      -- 
    cra_5008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2582_call_ack_0, ack => transmitEngineDaemon_CP_4738_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	84 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: 	43 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_Update/cca
      -- 
    cca_5013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2582_call_ack_1, ack => transmitEngineDaemon_CP_4738_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	56 
    -- CP-element group 68: 	59 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	76 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/barrier_stmt_2583_update_completed_
      -- 
    transmitEngineDaemon_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(67) & transmitEngineDaemon_CP_4738_elements(63) & transmitEngineDaemon_CP_4738_elements(56) & transmitEngineDaemon_CP_4738_elements(59);
      gj_transmitEngineDaemon_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Sample/req
      -- 
    req_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(69), ack => WPIPE_TX_ACTIVITY_LOGGER_2584_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(68) & transmitEngineDaemon_CP_4738_elements(71);
      gj_transmitEngineDaemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Sample/ack
      -- CP-element group 70: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Update/req
      -- 
    ack_5023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2584_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(70)); -- 
    req_5027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(70), ack => WPIPE_TX_ACTIVITY_LOGGER_2584_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	79 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2584_Update/ack
      -- 
    ack_5028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2584_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	84 
    -- CP-element group 72: 	52 
    -- CP-element group 72: 	59 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Sample/crr
      -- 
    crr_5036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(72), ack => call_stmt_2590_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(84) & transmitEngineDaemon_CP_4738_elements(52) & transmitEngineDaemon_CP_4738_elements(59);
      gj_transmitEngineDaemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Update/ccr
      -- 
    ccr_5041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(73), ack => call_stmt_2590_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_4738_elements(75);
      gj_transmitEngineDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	50 
    -- CP-element group 74: 	57 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Sample/cra
      -- 
    cra_5037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2590_call_ack_0, ack => transmitEngineDaemon_CP_4738_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	85 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	43 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2590_Update/cca
      -- CP-element group 75: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/ring_reenable_memory_space_0
      -- 
    cca_5042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2590_call_ack_1, ack => transmitEngineDaemon_CP_4738_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: 	25 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Sample/req
      -- 
    req_5050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(76), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(68) & transmitEngineDaemon_CP_4738_elements(25) & transmitEngineDaemon_CP_4738_elements(78);
      gj_transmitEngineDaemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	21 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Update/req
      -- 
    ack_5051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(77)); -- 
    req_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(77), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_Update/ack
      -- 
    ack_5056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/barrier_stmt_2594_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Sample/req
      -- 
    req_5065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(79), ack => WPIPE_TX_ACTIVITY_LOGGER_2595_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(71) & transmitEngineDaemon_CP_4738_elements(75) & transmitEngineDaemon_CP_4738_elements(78);
      gj_transmitEngineDaemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_update_start_
      -- CP-element group 80: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Update/req
      -- 
    ack_5066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2595_inst_ack_0, ack => transmitEngineDaemon_CP_4738_elements(80)); -- 
    req_5070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(80), ack => WPIPE_TX_ACTIVITY_LOGGER_2595_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	47 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/WPIPE_TX_ACTIVITY_LOGGER_2595_Update/ack
      -- 
    ack_5071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_TX_ACTIVITY_LOGGER_2595_inst_ack_1, ack => transmitEngineDaemon_CP_4738_elements(81)); -- 
    -- CP-element group 82:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	14 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	15 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_4738_elements(14), ack => transmitEngineDaemon_CP_4738_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	46 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	64 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2547_call_stmt_2582_delay
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_4738_elements(46), ack => transmitEngineDaemon_CP_4738_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	67 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	72 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/call_stmt_2582_call_stmt_2590_delay
      -- 
    -- Element group transmitEngineDaemon_CP_4738_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_4738_elements(67), ack => transmitEngineDaemon_CP_4738_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	17 
    -- CP-element group 85: 	18 
    -- CP-element group 85: 	75 
    -- CP-element group 85: 	81 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	11 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2509/do_while_stmt_2522/do_while_stmt_2522_loop_body/$exit
      -- 
    transmitEngineDaemon_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_4738_elements(17) & transmitEngineDaemon_CP_4738_elements(18) & transmitEngineDaemon_CP_4738_elements(75) & transmitEngineDaemon_CP_4738_elements(81);
      gj_transmitEngineDaemon_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	10 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_exit/$exit
      -- CP-element group 86: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_exit/ack
      -- 
    ack_5079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2522_branch_ack_0, ack => transmitEngineDaemon_CP_4738_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	10 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_taken/$exit
      -- CP-element group 87: 	 branch_block_stmt_2509/do_while_stmt_2522/loop_taken/ack
      -- 
    ack_5083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2522_branch_ack_1, ack => transmitEngineDaemon_CP_4738_elements(87)); -- 
    -- CP-element group 88:  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	8 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	4 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2509/do_while_stmt_2522/$exit
      -- 
    transmitEngineDaemon_CP_4738_elements(88) <= transmitEngineDaemon_CP_4738_elements(8);
    -- CP-element group 89:  merge  branch  transition  place  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	2 
    -- CP-element group 89: 	4 
    -- CP-element group 89: 	5 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	5 
    -- CP-element group 89: 	6 
    -- CP-element group 89:  members (49) 
      -- CP-element group 89: 	 branch_block_stmt_2509/merge_stmt_2510__exit__
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511__entry__
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_dead_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Sample/req
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Update/req
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/BITSEL_u32_u1_2514_inputs/RPIPE_S_CONTROL_REGISTER_2512/Update/ack
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/BITSEL_u32_u1_2514/SplitProtocol/Update/ca
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Update/cr
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/NOT_u1_u1_2515/SplitProtocol/Update/ca
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_eval_test/branch_req
      -- CP-element group 89: 	 branch_block_stmt_2509/NOT_u1_u1_2515_place
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_if_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/if_stmt_2511_else_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/merge_stmt_2510_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2509/merge_stmt_2510_PhiAck/$entry
      -- CP-element group 89: 	 branch_block_stmt_2509/merge_stmt_2510_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_2509/merge_stmt_2510_PhiAck/dummy
      -- 
    branch_req_4827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_4738_elements(89), ack => if_stmt_2511_branch_req_0); -- 
    transmitEngineDaemon_CP_4738_elements(89) <= OrReduce(transmitEngineDaemon_CP_4738_elements(2) & transmitEngineDaemon_CP_4738_elements(4) & transmitEngineDaemon_CP_4738_elements(5));
    transmitEngineDaemon_do_while_stmt_2522_terminator_5084: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_2522_terminator_5084", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_4738_elements(11),loop_continue => transmitEngineDaemon_CP_4738_elements(87),loop_terminate => transmitEngineDaemon_CP_4738_elements(86),loop_back => transmitEngineDaemon_CP_4738_elements(9),loop_exit => transmitEngineDaemon_CP_4738_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_2534_phi_seq_4913_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitEngineDaemon_CP_4738_elements(30);
      transmitEngineDaemon_CP_4738_elements(35)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitEngineDaemon_CP_4738_elements(35);
      transmitEngineDaemon_CP_4738_elements(36)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitEngineDaemon_CP_4738_elements(37);
      transmitEngineDaemon_CP_4738_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= transmitEngineDaemon_CP_4738_elements(32);
      transmitEngineDaemon_CP_4738_elements(39)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitEngineDaemon_CP_4738_elements(39);
      transmitEngineDaemon_CP_4738_elements(40)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitEngineDaemon_CP_4738_elements(41);
      transmitEngineDaemon_CP_4738_elements(33) <= phi_mux_reqs(1);
      phi_stmt_2534_phi_seq_4913 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2534_phi_seq_4913") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitEngineDaemon_CP_4738_elements(16), 
          phi_sample_ack => transmitEngineDaemon_CP_4738_elements(28), 
          phi_update_req => transmitEngineDaemon_CP_4738_elements(19), 
          phi_update_ack => transmitEngineDaemon_CP_4738_elements(29), 
          phi_mux_ack => transmitEngineDaemon_CP_4738_elements(34), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4856_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_4738_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_4738_elements(13);
        entry_tmerge_4856 : transition_merge -- 
          generic map(name => " entry_tmerge_4856")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_4738_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_2528_wire : std_logic_vector(7 downto 0);
    signal AND_u8_u8_2533_wire : std_logic_vector(7 downto 0);
    signal BITSEL_u32_u1_2514_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2601_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2466_2466_delayed_4_0_2564 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2515_wire : std_logic_vector(0 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_2526_wire : std_logic_vector(7 downto 0);
    signal RPIPE_S_CONTROL_REGISTER_2512_wire : std_logic_vector(31 downto 0);
    signal RPIPE_S_CONTROL_REGISTER_2599_wire : std_logic_vector(31 downto 0);
    signal RPIPE_S_NUMBER_OF_SERVERS_2529_wire : std_logic_vector(31 downto 0);
    signal R_FREEQUEUE_2578_wire_constant : std_logic_vector(1 downto 0);
    signal SUB_u32_u32_2531_wire : std_logic_vector(31 downto 0);
    signal init_flag_2534 : std_logic_vector(0 downto 0);
    signal konst_2507_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2513_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2527_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2530_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2550_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2559_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2579_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2585_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2596_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2600_wire_constant : std_logic_vector(31 downto 0);
    signal pkt_pointer_2477_delayed_4_0_2575 : std_logic_vector(63 downto 0);
    signal pkt_pointer_2547 : std_logic_vector(63 downto 0);
    signal push_pointer_back_to_free_Q_2569 : std_logic_vector(0 downto 0);
    signal push_status_2582 : std_logic_vector(0 downto 0);
    signal transmitted_flag_2556 : std_logic_vector(0 downto 0);
    signal tx_flag_2547 : std_logic_vector(0 downto 0);
    signal tx_q_index_2524 : std_logic_vector(7 downto 0);
    signal tx_tag_2520 : std_logic_vector(7 downto 0);
    signal type_cast_2532_wire : std_logic_vector(7 downto 0);
    signal type_cast_2537_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2539_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FREEQUEUE_2578_wire_constant <= "00";
    konst_2507_wire_constant <= "00000000";
    konst_2513_wire_constant <= "00000000000000000000000000000000";
    konst_2527_wire_constant <= "00000001";
    konst_2530_wire_constant <= "00000000000000000000000000000001";
    konst_2550_wire_constant <= "00000001";
    konst_2559_wire_constant <= "00000010";
    konst_2579_wire_constant <= "00000000";
    konst_2585_wire_constant <= "00000011";
    konst_2596_wire_constant <= "00000100";
    konst_2600_wire_constant <= "00000000000000000000000000000000";
    tx_tag_2520 <= "00000010";
    type_cast_2537_wire_constant <= "0";
    type_cast_2539_wire_constant <= "1";
    phi_stmt_2534: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2537_wire_constant & type_cast_2539_wire_constant;
      req <= phi_stmt_2534_req_0 & phi_stmt_2534_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2534",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2534_ack_0,
          idata => idata,
          odata => init_flag_2534,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2534
    W_pkt_pointer_2477_delayed_4_0_2573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_pointer_2477_delayed_4_0_2573_inst_req_0;
      W_pkt_pointer_2477_delayed_4_0_2573_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_pointer_2477_delayed_4_0_2573_inst_req_1;
      W_pkt_pointer_2477_delayed_4_0_2573_inst_ack_1<= rack(0);
      W_pkt_pointer_2477_delayed_4_0_2573_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_pointer_2477_delayed_4_0_2573_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_pointer_2547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_pointer_2477_delayed_4_0_2575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2524
    process(AND_u8_u8_2533_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := AND_u8_u8_2533_wire(7 downto 0);
      tx_q_index_2524 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2532_inst
    process(SUB_u32_u32_2531_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u32_u32_2531_wire(7 downto 0);
      type_cast_2532_wire <= tmp_var; -- 
    end process;
    do_while_stmt_2522_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_2601_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2522_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2522_branch_req_0,
          ack0 => do_while_stmt_2522_branch_ack_0,
          ack1 => do_while_stmt_2522_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2511_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2515_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2511_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2511_branch_req_0,
          ack0 => if_stmt_2511_branch_ack_0,
          ack1 => if_stmt_2511_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u8_u8_2528_inst
    ADD_u8_u8_2528_wire <= std_logic_vector(unsigned(RPIPE_LAST_READ_TX_QUEUE_INDEX_2526_wire) + unsigned(konst_2527_wire_constant));
    -- flow through binary operator AND_u1_u1_2568_inst
    push_pointer_back_to_free_Q_2569 <= (NOT_u1_u1_2466_2466_delayed_4_0_2564 and transmitted_flag_2556);
    -- shared split operator group (2) : AND_u8_u8_2533_inst 
    ApIntAnd_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u8_u8_2528_wire & type_cast_2532_wire;
      AND_u8_u8_2533_wire <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u8_u8_2533_inst_req_0;
      AND_u8_u8_2533_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u8_u8_2533_inst_req_1;
      AND_u8_u8_2533_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- flow through binary operator BITSEL_u32_u1_2514_inst
    process(RPIPE_S_CONTROL_REGISTER_2512_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_S_CONTROL_REGISTER_2512_wire, konst_2513_wire_constant, tmp_var);
      BITSEL_u32_u1_2514_wire <= tmp_var; --
    end process;
    -- flow through binary operator BITSEL_u32_u1_2601_inst
    process(RPIPE_S_CONTROL_REGISTER_2599_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_S_CONTROL_REGISTER_2599_wire, konst_2600_wire_constant, tmp_var);
      BITSEL_u32_u1_2601_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2515_inst
    process(BITSEL_u32_u1_2514_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_2514_wire, tmp_var);
      NOT_u1_u1_2515_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (6) : NOT_u1_u1_2563_inst 
    ApIntNot_group_6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tx_flag_2547;
      NOT_u1_u1_2466_2466_delayed_4_0_2564 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_2563_inst_req_0;
      NOT_u1_u1_2563_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_2563_inst_req_1;
      NOT_u1_u1_2563_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_6_gI: SplitGuardInterface generic map(name => "ApIntNot_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- flow through binary operator SUB_u32_u32_2531_inst
    SUB_u32_u32_2531_wire <= std_logic_vector(unsigned(RPIPE_S_NUMBER_OF_SERVERS_2529_wire) - unsigned(konst_2530_wire_constant));
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_2526_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- read from input-signal S_CONTROL_REGISTER
    RPIPE_S_CONTROL_REGISTER_2512_wire <= S_CONTROL_REGISTER;
    -- read from input-signal S_CONTROL_REGISTER
    RPIPE_S_CONTROL_REGISTER_2599_wire <= S_CONTROL_REGISTER;
    -- read from input-signal S_NUMBER_OF_SERVERS
    RPIPE_S_NUMBER_OF_SERVERS_2529_wire <= S_NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2506_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2507_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(15 downto 8),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2591_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_2524;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_TX_ACTIVITY_LOGGER_2584_inst WPIPE_TX_ACTIVITY_LOGGER_2558_inst WPIPE_TX_ACTIVITY_LOGGER_2549_inst WPIPE_TX_ACTIVITY_LOGGER_2595_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_TX_ACTIVITY_LOGGER_2584_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_TX_ACTIVITY_LOGGER_2558_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_TX_ACTIVITY_LOGGER_2549_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_TX_ACTIVITY_LOGGER_2595_inst_req_0;
      WPIPE_TX_ACTIVITY_LOGGER_2584_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_TX_ACTIVITY_LOGGER_2558_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_TX_ACTIVITY_LOGGER_2549_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_TX_ACTIVITY_LOGGER_2595_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_TX_ACTIVITY_LOGGER_2584_inst_req_1;
      update_req_unguarded(2) <= WPIPE_TX_ACTIVITY_LOGGER_2558_inst_req_1;
      update_req_unguarded(1) <= WPIPE_TX_ACTIVITY_LOGGER_2549_inst_req_1;
      update_req_unguarded(0) <= WPIPE_TX_ACTIVITY_LOGGER_2595_inst_req_1;
      WPIPE_TX_ACTIVITY_LOGGER_2584_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_TX_ACTIVITY_LOGGER_2558_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_TX_ACTIVITY_LOGGER_2549_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_TX_ACTIVITY_LOGGER_2595_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      data_in <= konst_2585_wire_constant & konst_2559_wire_constant & konst_2550_wire_constant & konst_2596_wire_constant;
      TX_ACTIVITY_LOGGER_write_2_gI: SplitGuardInterface generic map(name => "TX_ACTIVITY_LOGGER_write_2_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      TX_ACTIVITY_LOGGER_write_2: OutputPortRevised -- 
        generic map ( name => "TX_ACTIVITY_LOGGER", data_width => 8, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => TX_ACTIVITY_LOGGER_pipe_write_req(0),
          oack => TX_ACTIVITY_LOGGER_pipe_write_ack(0),
          odata => TX_ACTIVITY_LOGGER_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_2547_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2547_call_req_0;
      call_stmt_2547_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2547_call_req_1;
      call_stmt_2547_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_tag_2520 & tx_q_index_2524;
      pkt_pointer_2547 <= data_out(64 downto 1);
      tx_flag_2547 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 16,
        owidth => 16,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(15 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 65,
          owidth => 65,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(64 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2556_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2556_call_req_0;
      call_stmt_2556_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2556_call_req_1;
      call_stmt_2556_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not tx_flag_2547(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_tag_2520 & pkt_pointer_2547;
      transmitted_flag_2556 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(71 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2582_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(81 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2582_call_req_0;
      call_stmt_2582_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2582_call_req_1;
      call_stmt_2582_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_2569(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_tag_2520 & R_FREEQUEUE_2578_wire_constant & konst_2579_wire_constant & pkt_pointer_2477_delayed_4_0_2575;
      push_status_2582 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 82,
        owidth => 82,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(81 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2590_call 
    incrementNumberOfPacketsTransmitted_call_group_3: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2590_call_req_0;
      call_stmt_2590_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2590_call_req_1;
      call_stmt_2590_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_2569(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      incrementNumberOfPacketsTransmitted_call_group_3_gI: SplitGuardInterface generic map(name => "incrementNumberOfPacketsTransmitted_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => incrementNumberOfPacketsTransmitted_call_reqs(0),
          ackR => incrementNumberOfPacketsTransmitted_call_acks(0),
          tagR => incrementNumberOfPacketsTransmitted_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => incrementNumberOfPacketsTransmitted_return_acks(0), -- cross-over
          ackL => incrementNumberOfPacketsTransmitted_return_reqs(0), -- cross-over
          tagL => incrementNumberOfPacketsTransmitted_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    packet_pointer : in  std_logic_vector(63 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
    accessMemoryDword_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemoryDword_call_acks : in   std_logic_vector(1 downto 0);
    accessMemoryDword_call_data : out  std_logic_vector(401 downto 0);
    accessMemoryDword_call_tag  :  out  std_logic_vector(3 downto 0);
    accessMemoryDword_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemoryDword_return_acks : in   std_logic_vector(1 downto 0);
    accessMemoryDword_return_data : in   std_logic_vector(127 downto 0);
    accessMemoryDword_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal packet_pointer_buffer :  std_logic_vector(63 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_4465_start: Boolean;
  signal transmitPacket_CP_4465_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_2414_call_ack_1 : boolean;
  signal call_stmt_2414_call_req_1 : boolean;
  signal ncount_down_2462_2434_buf_req_1 : boolean;
  signal CONCAT_u65_u73_2456_inst_req_0 : boolean;
  signal CONCAT_u65_u73_2456_inst_ack_1 : boolean;
  signal CONCAT_u65_u73_2456_inst_ack_0 : boolean;
  signal ncount_down_2462_2434_buf_ack_1 : boolean;
  signal do_while_stmt_2427_branch_req_0 : boolean;
  signal CONCAT_u65_u73_2495_inst_ack_0 : boolean;
  signal W_last_offset_2475_inst_ack_1 : boolean;
  signal nmem_addr_offset_2467_2439_buf_req_1 : boolean;
  signal call_stmt_2449_call_req_0 : boolean;
  signal nmem_addr_offset_2467_2439_buf_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2450_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2450_inst_ack_0 : boolean;
  signal SUB_u11_u11_2433_inst_req_0 : boolean;
  signal call_stmt_2486_call_req_0 : boolean;
  signal SUB_u11_u11_2433_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2489_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2489_inst_req_1 : boolean;
  signal W_last_offset_2475_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2450_inst_req_1 : boolean;
  signal call_stmt_2486_call_req_1 : boolean;
  signal call_stmt_2486_call_ack_0 : boolean;
  signal CONCAT_u65_u73_2456_inst_req_1 : boolean;
  signal CONCAT_u65_u73_2495_inst_req_1 : boolean;
  signal phi_stmt_2435_req_1 : boolean;
  signal call_stmt_2486_call_ack_1 : boolean;
  signal EQ_u11_u1_2501_inst_ack_0 : boolean;
  signal SUB_u11_u11_2433_inst_req_1 : boolean;
  signal EQ_u11_u1_2501_inst_req_1 : boolean;
  signal EQ_u11_u1_2501_inst_req_0 : boolean;
  signal nmem_addr_offset_2467_2439_buf_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2450_inst_req_0 : boolean;
  signal EQ_u11_u1_2501_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2489_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2489_inst_ack_0 : boolean;
  signal nmem_addr_offset_2467_2439_buf_req_0 : boolean;
  signal call_stmt_2414_call_ack_0 : boolean;
  signal call_stmt_2414_call_req_0 : boolean;
  signal do_while_stmt_2427_branch_ack_1 : boolean;
  signal CONCAT_u65_u73_2495_inst_ack_1 : boolean;
  signal SUB_u11_u11_2433_inst_ack_1 : boolean;
  signal W_last_offset_2475_inst_req_1 : boolean;
  signal call_stmt_2449_call_ack_1 : boolean;
  signal ncount_down_2462_2434_buf_ack_0 : boolean;
  signal ncount_down_2462_2434_buf_req_0 : boolean;
  signal phi_stmt_2435_ack_0 : boolean;
  signal CONCAT_u65_u73_2495_inst_req_0 : boolean;
  signal phi_stmt_2429_ack_0 : boolean;
  signal do_while_stmt_2427_branch_ack_0 : boolean;
  signal call_stmt_2449_call_req_1 : boolean;
  signal phi_stmt_2435_req_0 : boolean;
  signal phi_stmt_2429_req_0 : boolean;
  signal call_stmt_2449_call_ack_0 : boolean;
  signal W_last_offset_2475_inst_ack_0 : boolean;
  signal phi_stmt_2429_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_4465_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_4465_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_4465_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_4465_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_4465: Block -- control-path 
    signal transmitPacket_CP_4465_elements: BooleanArray(82 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_4465_elements(0) <= transmitPacket_CP_4465_start;
    transmitPacket_CP_4465_symbol <= transmitPacket_CP_4465_elements(82);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Update/ccr
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_sample_start_
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_update_start_
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Update/$entry
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/$entry
      -- CP-element group 0: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Sample/crr
      -- CP-element group 0: 	 $entry
      -- 
    ccr_4483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(0), ack => call_stmt_2414_call_req_1); -- 
    crr_4478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(0), ack => call_stmt_2414_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_sample_completed_
      -- CP-element group 1: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Sample/cra
      -- CP-element group 1: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Sample/$exit
      -- 
    cra_4479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2414_call_ack_0, ack => transmitPacket_CP_4465_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_2426/branch_block_stmt_2426__entry__
      -- CP-element group 2: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2426/$entry
      -- CP-element group 2: 	 branch_block_stmt_2426/do_while_stmt_2427__entry__
      -- CP-element group 2: 	 assign_stmt_2403_to_assign_stmt_2422/call_stmt_2414_update_completed_
      -- CP-element group 2: 	 assign_stmt_2403_to_assign_stmt_2422/$exit
      -- 
    cca_4484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2414_call_ack_1, ack => transmitPacket_CP_4465_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	71 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3: 	73 
    -- CP-element group 3: 	75 
    -- CP-element group 3: 	77 
    -- CP-element group 3: 	81 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/$entry
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2426/do_while_stmt_2427__exit__
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502__entry__
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Sample/req
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Update/req
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_update_start_
      -- 
    req_4675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(3), ack => W_last_offset_2475_inst_req_0); -- 
    ccr_4694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(3), ack => call_stmt_2486_call_req_1); -- 
    cr_4708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(3), ack => CONCAT_u65_u73_2495_inst_req_1); -- 
    cr_4736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(3), ack => EQ_u11_u1_2501_inst_req_1); -- 
    req_4680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(3), ack => W_last_offset_2475_inst_req_1); -- 
    transmitPacket_CP_4465_elements(3) <= transmitPacket_CP_4465_elements(71);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_2426/do_while_stmt_2427/$entry
      -- CP-element group 4: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427__entry__
      -- 
    transmitPacket_CP_4465_elements(4) <= transmitPacket_CP_4465_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427__exit__
      -- 
    -- Element group transmitPacket_CP_4465_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_back
      -- 
    -- Element group transmitPacket_CP_4465_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	69 
    -- CP-element group 7: 	70 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_taken/$entry
      -- CP-element group 7: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_2426/do_while_stmt_2427/condition_done
      -- 
    transmitPacket_CP_4465_elements(7) <= transmitPacket_CP_4465_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	68 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_body_done
      -- 
    transmitPacket_CP_4465_elements(8) <= transmitPacket_CP_4465_elements(68);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	43 
    -- CP-element group 9: 	24 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/back_edge_to_loop_body
      -- 
    transmitPacket_CP_4465_elements(9) <= transmitPacket_CP_4465_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	45 
    -- CP-element group 10: 	26 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/first_time_through_loop_body
      -- 
    transmitPacket_CP_4465_elements(10) <= transmitPacket_CP_4465_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	39 
    -- CP-element group 11: 	40 
    -- CP-element group 11: 	67 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	19 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/$entry
      -- 
    -- Element group transmitPacket_CP_4465_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	67 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	23 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/condition_evaluated
      -- 
    condition_evaluated_4508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(12), ack => do_while_stmt_2427_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(67) & transmitPacket_CP_4465_elements(17) & transmitPacket_CP_4465_elements(23);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	39 
    -- CP-element group 13: 	18 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	20 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_sample_start__ps
      -- 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(39) & transmitPacket_CP_4465_elements(18) & transmitPacket_CP_4465_elements(17);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	41 
    -- CP-element group 14: 	21 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	68 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	18 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/aggregated_phi_sample_ack
      -- 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(41) & transmitPacket_CP_4465_elements(21);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	68 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group transmitPacket_CP_4465_elements(15) is a control-delay.
    cp_element_15_delay: control_delay_element  generic map(name => " 15_delay", delay_value => 1)  port map(req => transmitPacket_CP_4465_elements(14), ack => transmitPacket_CP_4465_elements(15), clk => clk, reset =>reset);
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	40 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/aggregated_phi_update_req
      -- CP-element group 16: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_update_start__ps
      -- 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(40) & transmitPacket_CP_4465_elements(19);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	42 
    -- CP-element group 17: 	23 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/aggregated_phi_update_ack
      -- 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(42) & transmitPacket_CP_4465_elements(23);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_sample_start_
      -- 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(11) & transmitPacket_CP_4465_elements(14);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	11 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_update_start_
      -- 
    transmitPacket_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(11) & transmitPacket_CP_4465_elements(23);
      gj_transmitPacket_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	13 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_sample_start__ps
      -- 
    transmitPacket_CP_4465_elements(20) <= transmitPacket_CP_4465_elements(13);
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	14 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_update_start__ps
      -- 
    transmitPacket_CP_4465_elements(22) <= transmitPacket_CP_4465_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: 	12 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	9 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_loopback_trigger
      -- 
    transmitPacket_CP_4465_elements(24) <= transmitPacket_CP_4465_elements(9);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_loopback_sample_req_ps
      -- CP-element group 25: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_loopback_sample_req
      -- 
    phi_stmt_2429_loopback_sample_req_4524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2429_loopback_sample_req_4524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(25), ack => phi_stmt_2429_req_1); -- 
    -- Element group transmitPacket_CP_4465_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	10 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_entry_trigger
      -- 
    transmitPacket_CP_4465_elements(26) <= transmitPacket_CP_4465_elements(10);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_entry_sample_req_ps
      -- CP-element group 27: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_entry_sample_req
      -- 
    phi_stmt_2429_entry_sample_req_4527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2429_entry_sample_req_4527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(27), ack => phi_stmt_2429_req_0); -- 
    -- Element group transmitPacket_CP_4465_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_phi_mux_ack_ps
      -- CP-element group 28: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2429_phi_mux_ack
      -- 
    phi_stmt_2429_phi_mux_ack_4530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2429_ack_0, ack => transmitPacket_CP_4465_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_update_start__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Sample/rr
      -- 
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(31), ack => SUB_u11_u11_2433_inst_req_0); -- 
    transmitPacket_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(29) & transmitPacket_CP_4465_elements(33);
      gj_transmitPacket_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Update/cr
      -- 
    cr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(32), ack => SUB_u11_u11_2433_inst_req_1); -- 
    transmitPacket_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(30) & transmitPacket_CP_4465_elements(34);
      gj_transmitPacket_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_sample_completed__ps
      -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u11_u11_2433_inst_ack_0, ack => transmitPacket_CP_4465_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/SUB_u11_u11_2433_Update/ca
      -- 
    ca_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u11_u11_2433_inst_ack_1, ack => transmitPacket_CP_4465_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_sample_start_
      -- 
    req_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(35), ack => ncount_down_2462_2434_buf_req_0); -- 
    -- Element group transmitPacket_CP_4465_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Update/req
      -- CP-element group 36: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_update_start_
      -- 
    req_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(36), ack => ncount_down_2462_2434_buf_req_1); -- 
    -- Element group transmitPacket_CP_4465_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_sample_completed_
      -- 
    ack_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_2462_2434_buf_ack_0, ack => transmitPacket_CP_4465_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Update/ack
      -- CP-element group 38: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_ncount_down_2434_update_completed__ps
      -- 
    ack_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_2462_2434_buf_ack_1, ack => transmitPacket_CP_4465_elements(38)); -- 
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	13 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_sample_start_
      -- 
    transmitPacket_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(11) & transmitPacket_CP_4465_elements(14);
      gj_transmitPacket_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	11 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: 	58 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	16 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_update_start_
      -- 
    transmitPacket_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(11) & transmitPacket_CP_4465_elements(42) & transmitPacket_CP_4465_elements(58);
      gj_transmitPacket_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	14 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	17 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	9 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_loopback_trigger
      -- 
    transmitPacket_CP_4465_elements(43) <= transmitPacket_CP_4465_elements(9);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_loopback_sample_req_ps
      -- 
    phi_stmt_2435_loopback_sample_req_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2435_loopback_sample_req_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(44), ack => phi_stmt_2435_req_1); -- 
    -- Element group transmitPacket_CP_4465_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_entry_trigger
      -- 
    transmitPacket_CP_4465_elements(45) <= transmitPacket_CP_4465_elements(10);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_entry_sample_req_ps
      -- CP-element group 46: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_entry_sample_req
      -- 
    phi_stmt_2435_entry_sample_req_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2435_entry_sample_req_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(46), ack => phi_stmt_2435_req_0); -- 
    -- Element group transmitPacket_CP_4465_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_phi_mux_ack_ps
      -- CP-element group 47: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/phi_stmt_2435_phi_mux_ack
      -- 
    phi_stmt_2435_phi_mux_ack_4584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2435_ack_0, ack => transmitPacket_CP_4465_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_update_start_
      -- CP-element group 49: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_update_start__ps
      -- 
    -- Element group transmitPacket_CP_4465_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_update_completed__ps
      -- 
    transmitPacket_CP_4465_elements(50) <= transmitPacket_CP_4465_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/type_cast_2438_update_completed_
      -- 
    -- Element group transmitPacket_CP_4465_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => transmitPacket_CP_4465_elements(49), ack => transmitPacket_CP_4465_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Sample/$entry
      -- 
    req_4605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(52), ack => nmem_addr_offset_2467_2439_buf_req_0); -- 
    -- Element group transmitPacket_CP_4465_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Update/req
      -- CP-element group 53: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_update_start_
      -- 
    req_4610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(53), ack => nmem_addr_offset_2467_2439_buf_req_1); -- 
    -- Element group transmitPacket_CP_4465_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Sample/$exit
      -- 
    ack_4606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_offset_2467_2439_buf_ack_0, ack => transmitPacket_CP_4465_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/R_nmem_addr_offset_2439_update_completed_
      -- 
    ack_4611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_offset_2467_2439_buf_ack_1, ack => transmitPacket_CP_4465_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Sample/crr
      -- CP-element group 56: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Sample/$entry
      -- 
    crr_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(56), ack => call_stmt_2449_call_req_0); -- 
    transmitPacket_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(42) & transmitPacket_CP_4465_elements(58);
      gj_transmitPacket_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	62 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Update/ccr
      -- CP-element group 57: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Update/$entry
      -- 
    ccr_4625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(57), ack => call_stmt_2449_call_req_1); -- 
    transmitPacket_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(59) & transmitPacket_CP_4465_elements(62);
      gj_transmitPacket_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	40 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Sample/cra
      -- 
    cra_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2449_call_ack_0, ack => transmitPacket_CP_4465_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Update/cca
      -- CP-element group 59: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/call_stmt_2449_Update/$exit
      -- 
    cca_4626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2449_call_ack_1, ack => transmitPacket_CP_4465_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_sample_start_
      -- 
    rr_4634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(60), ack => CONCAT_u65_u73_2456_inst_req_0); -- 
    transmitPacket_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(59) & transmitPacket_CP_4465_elements(62);
      gj_transmitPacket_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	65 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_update_start_
      -- CP-element group 61: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Update/cr
      -- 
    cr_4639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(61), ack => CONCAT_u65_u73_2456_inst_req_1); -- 
    transmitPacket_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(63) & transmitPacket_CP_4465_elements(65);
      gj_transmitPacket_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	57 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_sample_completed_
      -- 
    ra_4635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2456_inst_ack_0, ack => transmitPacket_CP_4465_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/CONCAT_u65_u73_2456_Update/$exit
      -- 
    ca_4640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2456_inst_ack_1, ack => transmitPacket_CP_4465_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_sample_start_
      -- 
    req_4648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(64), ack => WPIPE_nic_to_mac_transmit_pipe_2450_inst_req_0); -- 
    transmitPacket_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(63) & transmitPacket_CP_4465_elements(66);
      gj_transmitPacket_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	61 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Update/req
      -- CP-element group 65: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_sample_completed_
      -- 
    ack_4649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2450_inst_ack_0, ack => transmitPacket_CP_4465_elements(65)); -- 
    req_4653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(65), ack => WPIPE_nic_to_mac_transmit_pipe_2450_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/WPIPE_nic_to_mac_transmit_pipe_2450_update_completed_
      -- 
    ack_4654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2450_inst_ack_1, ack => transmitPacket_CP_4465_elements(66)); -- 
    -- CP-element group 67:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	11 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	12 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitPacket_CP_4465_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => transmitPacket_CP_4465_elements(11), ack => transmitPacket_CP_4465_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	14 
    -- CP-element group 68: 	15 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	8 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2426/do_while_stmt_2427/do_while_stmt_2427_loop_body/$exit
      -- 
    transmitPacket_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(66) & transmitPacket_CP_4465_elements(14) & transmitPacket_CP_4465_elements(15);
      gj_transmitPacket_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	7 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_exit/ack
      -- CP-element group 69: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_exit/$exit
      -- 
    ack_4659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2427_branch_ack_0, ack => transmitPacket_CP_4465_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	7 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_taken/ack
      -- CP-element group 70: 	 branch_block_stmt_2426/do_while_stmt_2427/loop_taken/$exit
      -- 
    ack_4663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2427_branch_ack_1, ack => transmitPacket_CP_4465_elements(70)); -- 
    -- CP-element group 71:  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	3 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2426/do_while_stmt_2427/$exit
      -- 
    transmitPacket_CP_4465_elements(71) <= transmitPacket_CP_4465_elements(5);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Sample/ack
      -- 
    ack_4676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_last_offset_2475_inst_ack_0, ack => transmitPacket_CP_4465_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	3 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	80 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Sample/crr
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/assign_stmt_2477_update_completed_
      -- 
    ack_4681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_last_offset_2475_inst_ack_1, ack => transmitPacket_CP_4465_elements(73)); -- 
    crr_4689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(73), ack => call_stmt_2486_call_req_0); -- 
    rr_4731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(73), ack => EQ_u11_u1_2501_inst_req_0); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Sample/cra
      -- CP-element group 74: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Sample/$exit
      -- 
    cra_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2486_call_ack_0, ack => transmitPacket_CP_4465_elements(74)); -- 
    -- CP-element group 75:  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	3 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (6) 
      -- CP-element group 75: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_Update/cca
      -- CP-element group 75: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/call_stmt_2486_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Sample/rr
      -- 
    cca_4695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2486_call_ack_1, ack => transmitPacket_CP_4465_elements(75)); -- 
    rr_4703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(75), ack => CONCAT_u65_u73_2495_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_sample_completed_
      -- 
    ra_4704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2495_inst_ack_0, ack => transmitPacket_CP_4465_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	3 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Sample/req
      -- CP-element group 77: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/CONCAT_u65_u73_2495_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Sample/$entry
      -- 
    ca_4709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2495_inst_ack_1, ack => transmitPacket_CP_4465_elements(77)); -- 
    req_4717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(77), ack => WPIPE_nic_to_mac_transmit_pipe_2489_inst_req_0); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Update/req
      -- CP-element group 78: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Sample/$exit
      -- 
    ack_4718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2489_inst_ack_0, ack => transmitPacket_CP_4465_elements(78)); -- 
    req_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_4465_elements(78), ack => WPIPE_nic_to_mac_transmit_pipe_2489_inst_req_1); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Update/ack
      -- CP-element group 79: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/WPIPE_nic_to_mac_transmit_pipe_2489_Update/$exit
      -- 
    ack_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2489_inst_ack_1, ack => transmitPacket_CP_4465_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	73 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_sample_completed_
      -- 
    ra_4732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u11_u1_2501_inst_ack_0, ack => transmitPacket_CP_4465_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	3 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/EQ_u11_u1_2501_Update/ca
      -- 
    ca_4737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u11_u1_2501_inst_ack_1, ack => transmitPacket_CP_4465_elements(81)); -- 
    -- CP-element group 82:  join  transition  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502/$exit
      -- CP-element group 82: 	 branch_block_stmt_2426/branch_block_stmt_2426__exit__
      -- CP-element group 82: 	 branch_block_stmt_2426/$exit
      -- CP-element group 82: 	 branch_block_stmt_2426/assign_stmt_2477_to_assign_stmt_2502__exit__
      -- CP-element group 82: 	 $exit
      -- 
    transmitPacket_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_4465_elements(79) & transmitPacket_CP_4465_elements(81);
      gj_transmitPacket_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_4465_elements(82), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_2427_terminator_4664: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_2427_terminator_4664", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_4465_elements(8),loop_continue => transmitPacket_CP_4465_elements(70),loop_terminate => transmitPacket_CP_4465_elements(69),loop_back => transmitPacket_CP_4465_elements(6),loop_exit => transmitPacket_CP_4465_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_2429_phi_seq_4568_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_4465_elements(26);
      transmitPacket_CP_4465_elements(29)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_4465_elements(33);
      transmitPacket_CP_4465_elements(30)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_4465_elements(34);
      transmitPacket_CP_4465_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_4465_elements(24);
      transmitPacket_CP_4465_elements(35)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_4465_elements(37);
      transmitPacket_CP_4465_elements(36)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_4465_elements(38);
      transmitPacket_CP_4465_elements(25) <= phi_mux_reqs(1);
      phi_stmt_2429_phi_seq_4568 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2429_phi_seq_4568") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_4465_elements(20), 
          phi_sample_ack => transmitPacket_CP_4465_elements(21), 
          phi_update_req => transmitPacket_CP_4465_elements(22), 
          phi_update_ack => transmitPacket_CP_4465_elements(23), 
          phi_mux_ack => transmitPacket_CP_4465_elements(28), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2435_phi_seq_4612_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_4465_elements(45);
      transmitPacket_CP_4465_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_4465_elements(48);
      transmitPacket_CP_4465_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_4465_elements(50);
      transmitPacket_CP_4465_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_4465_elements(43);
      transmitPacket_CP_4465_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_4465_elements(54);
      transmitPacket_CP_4465_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_4465_elements(55);
      transmitPacket_CP_4465_elements(44) <= phi_mux_reqs(1);
      phi_stmt_2435_phi_seq_4612 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2435_phi_seq_4612") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_4465_elements(13), 
          phi_sample_ack => transmitPacket_CP_4465_elements(41), 
          phi_update_req => transmitPacket_CP_4465_elements(16), 
          phi_update_ack => transmitPacket_CP_4465_elements(42), 
          phi_mux_ack => transmitPacket_CP_4465_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4509_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_4465_elements(9);
        preds(1)  <= transmitPacket_CP_4465_elements(10);
        entry_tmerge_4509 : transition_merge -- 
          generic map(name => " entry_tmerge_4509")
          port map (preds => preds, symbol_out => transmitPacket_CP_4465_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u65_2454_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_2493_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u65_u73_2456_wire : std_logic_vector(72 downto 0);
    signal CONCAT_u65_u73_2495_wire : std_logic_vector(72 downto 0);
    signal R_FULL_BYTE_MASK_2455_wire_constant : std_logic_vector(7 downto 0);
    signal R_READMEM_2408_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_2442_wire_constant : std_logic_vector(0 downto 0);
    signal R_READMEM_2479_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u11_u11_2433_wire : std_logic_vector(10 downto 0);
    signal control_data_2414 : std_logic_vector(63 downto 0);
    signal control_data_addr_2403 : std_logic_vector(63 downto 0);
    signal count_down_2429 : std_logic_vector(10 downto 0);
    signal data_2449 : std_logic_vector(63 downto 0);
    signal konst_2410_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2432_wire_constant : std_logic_vector(10 downto 0);
    signal konst_2460_wire_constant : std_logic_vector(10 downto 0);
    signal konst_2465_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2470_wire_constant : std_logic_vector(10 downto 0);
    signal last_offset_2477 : std_logic_vector(15 downto 0);
    signal last_tkeep_2422 : std_logic_vector(7 downto 0);
    signal last_word_2486 : std_logic_vector(63 downto 0);
    signal mem_addr_offset_2435 : std_logic_vector(15 downto 0);
    signal ncount_down_2462 : std_logic_vector(10 downto 0);
    signal ncount_down_2462_2434_buffered : std_logic_vector(10 downto 0);
    signal nmem_addr_offset_2467 : std_logic_vector(15 downto 0);
    signal nmem_addr_offset_2467_2439_buffered : std_logic_vector(15 downto 0);
    signal not_last_word_2472 : std_logic_vector(0 downto 0);
    signal packet_size_2418 : std_logic_vector(10 downto 0);
    signal type_cast_2412_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2438_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2445_wire : std_logic_vector(63 downto 0);
    signal type_cast_2447_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2452_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2482_wire : std_logic_vector(63 downto 0);
    signal type_cast_2484_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2491_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2500_wire : std_logic_vector(10 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_2455_wire_constant <= "11111111";
    R_READMEM_2408_wire_constant <= "1";
    R_READMEM_2442_wire_constant <= "1";
    R_READMEM_2479_wire_constant <= "1";
    konst_2410_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2432_wire_constant <= "00000010000";
    konst_2460_wire_constant <= "00000001000";
    konst_2465_wire_constant <= "0000000000001000";
    konst_2470_wire_constant <= "00000001000";
    type_cast_2412_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2438_wire_constant <= "0000000000011000";
    type_cast_2447_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2452_wire_constant <= "0";
    type_cast_2484_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2491_wire_constant <= "1";
    phi_stmt_2429: Block -- phi operator 
      signal idata: std_logic_vector(21 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SUB_u11_u11_2433_wire & ncount_down_2462_2434_buffered;
      req <= phi_stmt_2429_req_0 & phi_stmt_2429_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2429",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 11) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2429_ack_0,
          idata => idata,
          odata => count_down_2429,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2429
    phi_stmt_2435: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2438_wire_constant & nmem_addr_offset_2467_2439_buffered;
      req <= phi_stmt_2435_req_0 & phi_stmt_2435_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2435",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2435_ack_0,
          idata => idata,
          odata => mem_addr_offset_2435,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2435
    -- flow-through slice operator slice_2417_inst
    packet_size_2418 <= control_data_2414(18 downto 8);
    -- flow-through slice operator slice_2421_inst
    last_tkeep_2422 <= control_data_2414(7 downto 0);
    -- interlock W_control_data_addr_2401_inst
    process(packet_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := packet_pointer_buffer(63 downto 0);
      control_data_addr_2403 <= tmp_var; -- 
    end process;
    W_last_offset_2475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_last_offset_2475_inst_req_0;
      W_last_offset_2475_inst_ack_0<= wack(0);
      rreq(0) <= W_last_offset_2475_inst_req_1;
      W_last_offset_2475_inst_ack_1<= rack(0);
      W_last_offset_2475_inst : InterlockBuffer generic map ( -- 
        name => "W_last_offset_2475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_offset_2467,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => last_offset_2477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ncount_down_2462_2434_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_2462_2434_buf_req_0;
      ncount_down_2462_2434_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_2462_2434_buf_req_1;
      ncount_down_2462_2434_buf_ack_1<= rack(0);
      ncount_down_2462_2434_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_2462_2434_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 11,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_2462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_2462_2434_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmem_addr_offset_2467_2439_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_offset_2467_2439_buf_req_0;
      nmem_addr_offset_2467_2439_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_offset_2467_2439_buf_req_1;
      nmem_addr_offset_2467_2439_buf_ack_1<= rack(0);
      nmem_addr_offset_2467_2439_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_offset_2467_2439_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_offset_2467,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_offset_2467_2439_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2445_inst
    process(mem_addr_offset_2435) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mem_addr_offset_2435(15 downto 0);
      type_cast_2445_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2482_inst
    process(last_offset_2477) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := last_offset_2477(15 downto 0);
      type_cast_2482_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2500_inst
    process(last_offset_2477) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := last_offset_2477(10 downto 0);
      type_cast_2500_wire <= tmp_var; -- 
    end process;
    do_while_stmt_2427_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_2472;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2427_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2427_branch_req_0,
          ack0 => do_while_stmt_2427_branch_ack_0,
          ack1 => do_while_stmt_2427_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u16_u16_2466_inst
    nmem_addr_offset_2467 <= std_logic_vector(unsigned(mem_addr_offset_2435) + unsigned(konst_2465_wire_constant));
    -- flow through binary operator CONCAT_u1_u65_2454_inst
    process(type_cast_2452_wire_constant, data_2449) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2452_wire_constant, data_2449, tmp_var);
      CONCAT_u1_u65_2454_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u1_u65_2493_inst
    process(type_cast_2491_wire_constant, last_word_2486) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2491_wire_constant, last_word_2486, tmp_var);
      CONCAT_u1_u65_2493_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : CONCAT_u65_u73_2456_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_2454_wire;
      CONCAT_u65_u73_2456_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_2456_inst_req_0;
      CONCAT_u65_u73_2456_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_2456_inst_req_1;
      CONCAT_u65_u73_2456_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : CONCAT_u65_u73_2495_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_2493_wire & last_tkeep_2422;
      CONCAT_u65_u73_2495_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_2495_inst_req_0;
      CONCAT_u65_u73_2495_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_2495_inst_req_1;
      CONCAT_u65_u73_2495_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : EQ_u11_u1_2501_inst 
    ApIntEq_group_5: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_2418 & type_cast_2500_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u11_u1_2501_inst_req_0;
      EQ_u11_u1_2501_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u11_u1_2501_inst_req_1;
      EQ_u11_u1_2501_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_5_gI: SplitGuardInterface generic map(name => "ApIntEq_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : SUB_u11_u11_2433_inst 
    ApIntSub_group_6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_2418;
      SUB_u11_u11_2433_wire <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u11_u11_2433_inst_req_0;
      SUB_u11_u11_2433_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u11_u11_2433_inst_req_1;
      SUB_u11_u11_2433_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_6_gI: SplitGuardInterface generic map(name => "ApIntSub_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000010000",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- flow through binary operator SUB_u11_u11_2461_inst
    ncount_down_2462 <= std_logic_vector(unsigned(count_down_2429) - unsigned(konst_2460_wire_constant));
    -- flow through binary operator UGT_u11_u1_2471_inst
    process(ncount_down_2462) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_2462, konst_2470_wire_constant, tmp_var);
      not_last_word_2472 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_2450_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2450_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_2450_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2450_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_2450_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_2456_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(1),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(1),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 73),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_to_mac_transmit_pipe_2489_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2489_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_2489_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2489_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_2489_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_2495_wire;
      nic_to_mac_transmit_pipe_write_1_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2486_call call_stmt_2414_call 
    accessMemoryDword_call_group_0: Block -- 
      signal data_in: std_logic_vector(401 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2486_call_req_0;
      reqL_unguarded(0) <= call_stmt_2414_call_req_0;
      call_stmt_2486_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2414_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2486_call_req_1;
      reqR_unguarded(0) <= call_stmt_2414_call_req_1;
      call_stmt_2486_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2414_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemoryDword_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemoryDword_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemoryDword_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemoryDword_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemoryDword_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_2479_wire_constant & control_data_addr_2403 & type_cast_2482_wire & type_cast_2484_wire_constant & tag_buffer & R_READMEM_2408_wire_constant & control_data_addr_2403 & konst_2410_wire_constant & type_cast_2412_wire_constant;
      last_word_2486 <= data_out(127 downto 64);
      control_data_2414 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 402,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(1),
          ackR => accessMemoryDword_call_acks(1),
          dataR => accessMemoryDword_call_data(401 downto 201),
          tagR => accessMemoryDword_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(1), -- cross-over
          ackL => accessMemoryDword_return_reqs(1), -- cross-over
          dataL => accessMemoryDword_return_data(127 downto 64),
          tagL => accessMemoryDword_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2449_call 
    accessMemoryDword_call_group_1: Block -- 
      signal data_in: std_logic_vector(200 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 38);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2449_call_req_0;
      call_stmt_2449_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2449_call_req_1;
      call_stmt_2449_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDword_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tag_buffer & R_READMEM_2442_wire_constant & control_data_addr_2403 & type_cast_2445_wire & type_cast_2447_wire_constant;
      data_2449 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 201,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(0),
          ackR => accessMemoryDword_call_acks(0),
          dataR => accessMemoryDword_call_data(200 downto 0),
          tagR => accessMemoryDword_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(0), -- cross-over
          ackL => accessMemoryDword_return_reqs(0), -- cross-over
          dataL => accessMemoryDword_return_data(63 downto 0),
          tagL => accessMemoryDword_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    base_buffer_pointer : in  std_logic_vector(63 downto 0);
    max_addr_offset : in  std_logic_vector(15 downto 0);
    packet_size : in  std_logic_vector(10 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
    accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
    accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 107)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal base_buffer_pointer_buffer :  std_logic_vector(63 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal max_addr_offset_buffer :  std_logic_vector(15 downto 0);
  signal max_addr_offset_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(10 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_2230_start: Boolean;
  signal writeControlInformationToMem_CP_2230_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1512_call_ack_1 : boolean;
  signal call_stmt_1512_call_req_1 : boolean;
  signal call_stmt_1512_call_ack_0 : boolean;
  signal call_stmt_1512_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 107) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(87 downto 72) <= max_addr_offset;
  max_addr_offset_buffer <= in_buffer_data_out(87 downto 72);
  in_buffer_data_in(98 downto 88) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(98 downto 88);
  in_buffer_data_in(106 downto 99) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(106 downto 99);
  in_buffer_data_in(tag_length + 106 downto 107) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 106 downto 107);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_2230_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_2230_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_2230_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_2230_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_2230: Block -- control-path 
    signal writeControlInformationToMem_CP_2230_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_2230_elements(0) <= writeControlInformationToMem_CP_2230_start;
    writeControlInformationToMem_CP_2230_symbol <= writeControlInformationToMem_CP_2230_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_sample_start_
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_update_start_
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1497_to_call_stmt_1512/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_2230_elements(0), ack => call_stmt_1512_call_req_0); -- 
    ccr_2248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_2230_elements(0), ack => call_stmt_1512_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Sample/cra
      -- 
    cra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1512_call_ack_0, ack => writeControlInformationToMem_CP_2230_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_update_completed_
      -- CP-element group 2: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Update/cca
      -- CP-element group 2: 	 assign_stmt_1497_to_call_stmt_1512/call_stmt_1512_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1497_to_call_stmt_1512/$exit
      -- CP-element group 2: 	 $exit
      -- 
    cca_2249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1512_call_ack_1, ack => writeControlInformationToMem_CP_2230_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u11_u19_1495_wire : std_logic_vector(18 downto 0);
    signal CONCAT_u16_u45_1492_wire : std_logic_vector(44 downto 0);
    signal R_WRITEMEM_1507_wire_constant : std_logic_vector(0 downto 0);
    signal SHL_u8_u8_1501_wire : std_logic_vector(7 downto 0);
    signal control_data_1497 : std_logic_vector(63 downto 0);
    signal ctrlInfoTag_1505 : std_logic_vector(7 downto 0);
    signal ignore_return_1512 : std_logic_vector(63 downto 0);
    signal konst_1500_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1509_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1491_wire_constant : std_logic_vector(28 downto 0);
    signal type_cast_1503_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_WRITEMEM_1507_wire_constant <= "0";
    konst_1500_wire_constant <= "00000010";
    konst_1509_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1491_wire_constant <= "00000000000000000000000000000";
    type_cast_1503_wire_constant <= "00000011";
    -- flow through binary operator CONCAT_u11_u19_1495_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(18 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u11_u19_1495_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u16_u45_1492_inst
    process(max_addr_offset_buffer) -- 
      variable tmp_var : std_logic_vector(44 downto 0); -- 
    begin -- 
      ApConcat_proc(max_addr_offset_buffer, type_cast_1491_wire_constant, tmp_var);
      CONCAT_u16_u45_1492_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u45_u64_1496_inst
    process(CONCAT_u16_u45_1492_wire, CONCAT_u11_u19_1495_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u45_1492_wire, CONCAT_u11_u19_1495_wire, tmp_var);
      control_data_1497 <= tmp_var; --
    end process;
    -- flow through binary operator OR_u8_u8_1504_inst
    ctrlInfoTag_1505 <= (SHL_u8_u8_1501_wire or type_cast_1503_wire_constant);
    -- flow through binary operator SHL_u8_u8_1501_inst
    process(tag_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tag_buffer, konst_1500_wire_constant, tmp_var);
      SHL_u8_u8_1501_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1512_call 
    accessMemoryDword_call_group_0: Block -- 
      signal data_in: std_logic_vector(200 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1512_call_req_0;
      call_stmt_1512_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1512_call_req_1;
      call_stmt_1512_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDword_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ctrlInfoTag_1505 & R_WRITEMEM_1507_wire_constant & base_buffer_pointer_buffer & konst_1509_wire_constant & control_data_1497;
      ignore_return_1512 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 201,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(0),
          ackR => accessMemoryDword_call_acks(0),
          dataR => accessMemoryDword_call_data(200 downto 0),
          tagR => accessMemoryDword_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(0), -- cross-over
          ackL => accessMemoryDword_return_reqs(0), -- cross-over
          dataL => accessMemoryDword_return_data(63 downto 0),
          tagL => accessMemoryDword_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    buf_pointer : in  std_logic_vector(63 downto 0);
    addr_offset : out  std_logic_vector(15 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
    accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
    accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(63 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal addr_offset_buffer :  std_logic_vector(15 downto 0);
  signal addr_offset_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_1925_start: Boolean;
  signal writeEthernetHeaderToMem_CP_1925_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal naddr_offset_1385_1355_buf_ack_0 : boolean;
  signal do_while_stmt_1349_branch_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_1364_inst_req_0 : boolean;
  signal phi_stmt_1356_req_0 : boolean;
  signal call_stmt_1380_call_ack_1 : boolean;
  signal do_while_stmt_1349_branch_ack_1 : boolean;
  signal phi_stmt_1351_req_0 : boolean;
  signal phi_stmt_1356_ack_0 : boolean;
  signal call_stmt_1380_call_req_1 : boolean;
  signal phi_stmt_1351_req_1 : boolean;
  signal naddr_offset_1385_1355_buf_req_0 : boolean;
  signal RPIPE_nic_rx_to_header_1364_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_1364_inst_ack_1 : boolean;
  signal type_cast_1372_inst_req_0 : boolean;
  signal type_cast_1372_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_1364_inst_req_1 : boolean;
  signal phi_stmt_1356_req_1 : boolean;
  signal call_stmt_1380_call_ack_0 : boolean;
  signal call_stmt_1380_call_req_0 : boolean;
  signal type_cast_1372_inst_ack_1 : boolean;
  signal type_cast_1372_inst_req_1 : boolean;
  signal phi_stmt_1351_ack_0 : boolean;
  signal naddr_offset_1385_1355_buf_ack_1 : boolean;
  signal naddr_offset_1385_1355_buf_req_1 : boolean;
  signal do_while_stmt_1349_branch_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(71 downto 8) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 8);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_1925_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= addr_offset_buffer;
  addr_offset <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1925_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1925_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1925_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_1925: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_1925_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_1925_elements(0) <= writeEthernetHeaderToMem_CP_1925_start;
    writeEthernetHeaderToMem_CP_1925_symbol <= writeEthernetHeaderToMem_CP_1925_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1340/assign_stmt_1348/$exit
      -- CP-element group 0: 	 branch_block_stmt_1340/assign_stmt_1348/$entry
      -- CP-element group 0: 	 branch_block_stmt_1340/do_while_stmt_1349__entry__
      -- CP-element group 0: 	 branch_block_stmt_1340/assign_stmt_1348__exit__
      -- CP-element group 0: 	 branch_block_stmt_1340/$entry
      -- CP-element group 0: 	 branch_block_stmt_1340/assign_stmt_1348__entry__
      -- CP-element group 0: 	 branch_block_stmt_1340/branch_block_stmt_1340__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	68 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1340/do_while_stmt_1349__exit__
      -- CP-element group 1: 	 branch_block_stmt_1340/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1340/branch_block_stmt_1340__exit__
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(1) <= writeEthernetHeaderToMem_CP_1925_elements(68);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1340/do_while_stmt_1349/$entry
      -- CP-element group 2: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349__entry__
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(2) <= writeEthernetHeaderToMem_CP_1925_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	68 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349__exit__
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_back
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	66 
    -- CP-element group 5: 	67 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1340/do_while_stmt_1349/condition_done
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(5) <= writeEthernetHeaderToMem_CP_1925_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	65 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_body_done
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(6) <= writeEthernetHeaderToMem_CP_1925_elements(65);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	39 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/back_edge_to_loop_body
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(7) <= writeEthernetHeaderToMem_CP_1925_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8: 	41 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/first_time_through_loop_body
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(8) <= writeEthernetHeaderToMem_CP_1925_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	64 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	52 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1362_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/loop_body_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	64 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/condition_evaluated
      -- 
    condition_evaluated_1954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(10), ack => do_while_stmt_1349_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(64) & writeEthernetHeaderToMem_CP_1925_elements(15);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	33 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	53 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_sample_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(9) & writeEthernetHeaderToMem_CP_1925_elements(16) & writeEthernetHeaderToMem_CP_1925_elements(33) & writeEthernetHeaderToMem_CP_1925_elements(15);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	55 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: 	13 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1362_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_sample_completed_
      -- 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(18) & writeEthernetHeaderToMem_CP_1925_elements(36) & writeEthernetHeaderToMem_CP_1925_elements(55);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	65 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1925_elements(12), ack => writeEthernetHeaderToMem_CP_1925_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	34 
    -- CP-element group 14: 	52 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	54 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_update_start__ps
      -- CP-element group 14: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/aggregated_phi_update_req
      -- 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(17) & writeEthernetHeaderToMem_CP_1925_elements(34) & writeEthernetHeaderToMem_CP_1925_elements(52);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	56 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/aggregated_phi_update_ack
      -- 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(19) & writeEthernetHeaderToMem_CP_1925_elements(38) & writeEthernetHeaderToMem_CP_1925_elements(56);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(9) & writeEthernetHeaderToMem_CP_1925_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	58 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(9) & writeEthernetHeaderToMem_CP_1925_elements(58);
      gj_writeEthernetHeaderToMem_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	58 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_update_completed__ps
      -- CP-element group 19: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_update_completed_
      -- 
    rr_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(19), ack => type_cast_1372_inst_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(20) <= writeEthernetHeaderToMem_CP_1925_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_loopback_sample_req
      -- CP-element group 21: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_loopback_sample_req_ps
      -- 
    phi_stmt_1351_loopback_sample_req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1351_loopback_sample_req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(21), ack => phi_stmt_1351_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(22) <= writeEthernetHeaderToMem_CP_1925_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_entry_sample_req_ps
      -- CP-element group 23: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_entry_sample_req
      -- 
    phi_stmt_1351_entry_sample_req_1973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1351_entry_sample_req_1973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(23), ack => phi_stmt_1351_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_phi_mux_ack_ps
      -- CP-element group 24: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1351_phi_mux_ack
      -- 
    phi_stmt_1351_phi_mux_ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1351_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(27) <= writeEthernetHeaderToMem_CP_1925_elements(28);
    -- CP-element group 28:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	27 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1354_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1925_elements(26), ack => writeEthernetHeaderToMem_CP_1925_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_sample_start_
      -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(29), ack => naddr_offset_1385_1355_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Update/req
      -- 
    req_2002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(30), ack => naddr_offset_1385_1355_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_sample_completed_
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => naddr_offset_1385_1355_buf_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(31)); -- 
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/R_naddr_offset_1355_Update/ack
      -- 
    ack_2003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => naddr_offset_1385_1355_buf_ack_1, ack => writeEthernetHeaderToMem_CP_1925_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	12 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	11 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(9) & writeEthernetHeaderToMem_CP_1925_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	38 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	14 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(9) & writeEthernetHeaderToMem_CP_1925_elements(38);
      gj_writeEthernetHeaderToMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_sample_start__ps
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(35) <= writeEthernetHeaderToMem_CP_1925_elements(11);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	12 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(36) is bound as output of CP function.
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_update_start__ps
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(37) <= writeEthernetHeaderToMem_CP_1925_elements(14);
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	34 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	7 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(39) <= writeEthernetHeaderToMem_CP_1925_elements(7);
    -- CP-element group 40:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_loopback_sample_req_ps
      -- CP-element group 40: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_loopback_sample_req
      -- 
    phi_stmt_1356_loopback_sample_req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1356_loopback_sample_req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(40), ack => phi_stmt_1356_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	8 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(41) <= writeEthernetHeaderToMem_CP_1925_elements(8);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_entry_sample_req_ps
      -- CP-element group 42: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_entry_sample_req
      -- 
    phi_stmt_1356_entry_sample_req_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1356_entry_sample_req_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(42), ack => phi_stmt_1356_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_phi_mux_ack_ps
      -- CP-element group 43: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1356_phi_mux_ack
      -- 
    phi_stmt_1356_phi_mux_ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1356_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_sample_start__ps
      -- CP-element group 44: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_sample_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_sample_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_update_start__ps
      -- CP-element group 45: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_update_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(46) <= writeEthernetHeaderToMem_CP_1925_elements(47);
    -- CP-element group 47:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	46 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1359_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(47) is a control-delay.
    cp_element_47_delay: control_delay_element  generic map(name => " 47_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1925_elements(45), ack => writeEthernetHeaderToMem_CP_1925_elements(47), clk => clk, reset =>reset);
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_update_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(50) <= writeEthernetHeaderToMem_CP_1925_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1361_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1925_elements(49), ack => writeEthernetHeaderToMem_CP_1925_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	62 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	14 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1362_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(9) & writeEthernetHeaderToMem_CP_1925_elements(62);
      gj_writeEthernetHeaderToMem_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Sample/$entry
      -- 
    rr_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(53), ack => RPIPE_nic_rx_to_header_1364_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(11) & writeEthernetHeaderToMem_CP_1925_elements(56);
      gj_writeEthernetHeaderToMem_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	14 
    -- CP-element group 54: 	55 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Update/cr
      -- 
    cr_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(54), ack => RPIPE_nic_rx_to_header_1364_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(14) & writeEthernetHeaderToMem_CP_1925_elements(55);
      gj_writeEthernetHeaderToMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: 	54 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Sample/$exit
      -- 
    ra_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_1364_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	15 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/phi_stmt_1362_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/RPIPE_nic_rx_to_header_1364_Update/$exit
      -- 
    ca_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_1364_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1925_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	62 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Update/cr
      -- 
    cr_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(57), ack => type_cast_1372_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_1925_elements(62);
      gj_writeEthernetHeaderToMem_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	19 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	17 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Sample/ra
      -- 
    ra_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1372_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/type_cast_1372_Update/ca
      -- 
    ca_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1372_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1925_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: 	56 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Sample/crr
      -- CP-element group 60: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Sample/$entry
      -- 
    crr_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(60), ack => call_stmt_1380_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(59) & writeEthernetHeaderToMem_CP_1925_elements(56);
      gj_writeEthernetHeaderToMem_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Update/ccr
      -- CP-element group 61: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_update_start_
      -- 
    ccr_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1925_elements(61), ack => call_stmt_1380_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_1925_elements(63);
      gj_writeEthernetHeaderToMem_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	57 
    -- CP-element group 62: 	52 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Sample/cra
      -- CP-element group 62: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Sample/$exit
      -- 
    cra_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1380_call_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Update/cca
      -- CP-element group 63: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/call_stmt_1380_update_completed_
      -- 
    cca_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1380_call_ack_1, ack => writeEthernetHeaderToMem_CP_1925_elements(63)); -- 
    -- CP-element group 64:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	9 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	10 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1925_elements(64) is a control-delay.
    cp_element_64_delay: control_delay_element  generic map(name => " 64_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1925_elements(9), ack => writeEthernetHeaderToMem_CP_1925_elements(64), clk => clk, reset =>reset);
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	13 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	6 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1340/do_while_stmt_1349/do_while_stmt_1349_loop_body/$exit
      -- 
    writeEthernetHeaderToMem_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1925_elements(63) & writeEthernetHeaderToMem_CP_1925_elements(12) & writeEthernetHeaderToMem_CP_1925_elements(13);
      gj_writeEthernetHeaderToMem_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	5 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_exit/$exit
      -- CP-element group 66: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_exit/ack
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1349_branch_ack_0, ack => writeEthernetHeaderToMem_CP_1925_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	5 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_taken/$exit
      -- CP-element group 67: 	 branch_block_stmt_1340/do_while_stmt_1349/loop_taken/ack
      -- 
    ack_2093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1349_branch_ack_1, ack => writeEthernetHeaderToMem_CP_1925_elements(67)); -- 
    -- CP-element group 68:  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	3 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	1 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1340/do_while_stmt_1349/$exit
      -- 
    writeEthernetHeaderToMem_CP_1925_elements(68) <= writeEthernetHeaderToMem_CP_1925_elements(3);
    writeEthernetHeaderToMem_do_while_stmt_1349_terminator_2094: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_1349_terminator_2094", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_1925_elements(6),loop_continue => writeEthernetHeaderToMem_CP_1925_elements(67),loop_terminate => writeEthernetHeaderToMem_CP_1925_elements(66),loop_back => writeEthernetHeaderToMem_CP_1925_elements(4),loop_exit => writeEthernetHeaderToMem_CP_1925_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1351_phi_seq_2004_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_1925_elements(22);
      writeEthernetHeaderToMem_CP_1925_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_1925_elements(25);
      writeEthernetHeaderToMem_CP_1925_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_1925_elements(27);
      writeEthernetHeaderToMem_CP_1925_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_1925_elements(20);
      writeEthernetHeaderToMem_CP_1925_elements(29)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_1925_elements(31);
      writeEthernetHeaderToMem_CP_1925_elements(30)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_1925_elements(32);
      writeEthernetHeaderToMem_CP_1925_elements(21) <= phi_mux_reqs(1);
      phi_stmt_1351_phi_seq_2004 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1351_phi_seq_2004") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_1925_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_1925_elements(18), 
          phi_update_req => writeEthernetHeaderToMem_CP_1925_elements(14), 
          phi_update_ack => writeEthernetHeaderToMem_CP_1925_elements(19), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_1925_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1356_phi_seq_2038_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_1925_elements(41);
      writeEthernetHeaderToMem_CP_1925_elements(44)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_1925_elements(44);
      writeEthernetHeaderToMem_CP_1925_elements(45)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_1925_elements(46);
      writeEthernetHeaderToMem_CP_1925_elements(42) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_1925_elements(39);
      writeEthernetHeaderToMem_CP_1925_elements(48)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_1925_elements(48);
      writeEthernetHeaderToMem_CP_1925_elements(49)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_1925_elements(50);
      writeEthernetHeaderToMem_CP_1925_elements(40) <= phi_mux_reqs(1);
      phi_stmt_1356_phi_seq_2038 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1356_phi_seq_2038") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_1925_elements(35), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_1925_elements(36), 
          phi_update_req => writeEthernetHeaderToMem_CP_1925_elements(37), 
          phi_update_ack => writeEthernetHeaderToMem_CP_1925_elements(38), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_1925_elements(43), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1955_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_1925_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_1925_elements(8);
        entry_tmerge_1955 : transition_merge -- 
          generic map(name => " entry_tmerge_1955")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1925_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_nic_rx_to_header_1364_wire : std_logic_vector(72 downto 0);
    signal R_WRITEMEM_1375_wire_constant : std_logic_vector(0 downto 0);
    signal SHL_u8_u8_1344_wire : std_logic_vector(7 downto 0);
    signal ethHeaderTag_1348 : std_logic_vector(7 downto 0);
    signal ethernet_header_1362 : std_logic_vector(72 downto 0);
    signal first_time_1356 : std_logic_vector(0 downto 0);
    signal ignore_return_1380 : std_logic_vector(63 downto 0);
    signal konst_1343_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1383_wire_constant : std_logic_vector(15 downto 0);
    signal naddr_offset_1385 : std_logic_vector(15 downto 0);
    signal naddr_offset_1385_1355_buffered : std_logic_vector(15 downto 0);
    signal type_cast_1307_1307_delayed_1_0_1373 : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1354_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1361_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_1369 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    R_WRITEMEM_1375_wire_constant <= "0";
    konst_1343_wire_constant <= "00000010";
    konst_1383_wire_constant <= "0000000000001000";
    type_cast_1346_wire_constant <= "00000001";
    type_cast_1354_wire_constant <= "0000000000001000";
    type_cast_1359_wire_constant <= "1";
    type_cast_1361_wire_constant <= "0";
    phi_stmt_1351: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1354_wire_constant & naddr_offset_1385_1355_buffered;
      req <= phi_stmt_1351_req_0 & phi_stmt_1351_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1351",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1351_ack_0,
          idata => idata,
          odata => addr_offset_buffer,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1351
    phi_stmt_1356: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1359_wire_constant & type_cast_1361_wire_constant;
      req <= phi_stmt_1356_req_0 & phi_stmt_1356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1356",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1356_ack_0,
          idata => idata,
          odata => first_time_1356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1356
    -- flow-through slice operator slice_1368_inst
    wdata_1369 <= ethernet_header_1362(71 downto 8);
    naddr_offset_1385_1355_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= naddr_offset_1385_1355_buf_req_0;
      naddr_offset_1385_1355_buf_ack_0<= wack(0);
      rreq(0) <= naddr_offset_1385_1355_buf_req_1;
      naddr_offset_1385_1355_buf_ack_1<= rack(0);
      naddr_offset_1385_1355_buf : InterlockBuffer generic map ( -- 
        name => "naddr_offset_1385_1355_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => naddr_offset_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => naddr_offset_1385_1355_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1362
    process(RPIPE_nic_rx_to_header_1364_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_1364_wire(72 downto 0);
      ethernet_header_1362 <= tmp_var; -- 
    end process;
    type_cast_1372_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1372_inst_req_0;
      type_cast_1372_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1372_inst_req_1;
      type_cast_1372_inst_ack_1<= rack(0);
      type_cast_1372_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1372_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => addr_offset_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1307_1307_delayed_1_0_1373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1349_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= first_time_1356;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1349_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1349_branch_req_0,
          ack0 => do_while_stmt_1349_branch_ack_0,
          ack1 => do_while_stmt_1349_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u16_u16_1384_inst
    naddr_offset_1385 <= std_logic_vector(unsigned(addr_offset_buffer) + unsigned(konst_1383_wire_constant));
    -- flow through binary operator OR_u8_u8_1347_inst
    ethHeaderTag_1348 <= (SHL_u8_u8_1344_wire or type_cast_1346_wire_constant);
    -- flow through binary operator SHL_u8_u8_1344_inst
    process(tag_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tag_buffer, konst_1343_wire_constant, tmp_var);
      SHL_u8_u8_1344_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_1364_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_1364_inst_req_0;
      RPIPE_nic_rx_to_header_1364_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_1364_inst_req_1;
      RPIPE_nic_rx_to_header_1364_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_1364_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1380_call 
    accessMemoryDword_call_group_0: Block -- 
      signal data_in: std_logic_vector(200 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 38);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1380_call_req_0;
      call_stmt_1380_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1380_call_req_1;
      call_stmt_1380_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDword_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ethHeaderTag_1348 & R_WRITEMEM_1375_wire_constant & buf_pointer_buffer & type_cast_1307_1307_delayed_1_0_1373 & wdata_1369;
      ignore_return_1380 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 201,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(0),
          ackR => accessMemoryDword_call_acks(0),
          dataR => accessMemoryDword_call_data(200 downto 0),
          tagR => accessMemoryDword_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(0), -- cross-over
          ackL => accessMemoryDword_return_reqs(0), -- cross-over
          dataL => accessMemoryDword_return_data(63 downto 0),
          tagL => accessMemoryDword_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    tag : in  std_logic_vector(7 downto 0);
    max_addr_offset : in  std_logic_vector(15 downto 0);
    base_buf_pointer : in  std_logic_vector(63 downto 0);
    addr_offset : in  std_logic_vector(15 downto 0);
    packet_size_11 : out  std_logic_vector(10 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
    accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
    accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
    accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 20)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal tag_buffer :  std_logic_vector(7 downto 0);
  signal tag_update_enable: Boolean;
  signal max_addr_offset_buffer :  std_logic_vector(15 downto 0);
  signal max_addr_offset_update_enable: Boolean;
  signal base_buf_pointer_buffer :  std_logic_vector(63 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal addr_offset_buffer :  std_logic_vector(15 downto 0);
  signal addr_offset_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_11_buffer :  std_logic_vector(10 downto 0);
  signal packet_size_11_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_2095_start: Boolean;
  signal writePayloadToMem_CP_2095_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_1408_branch_req_0 : boolean;
  signal phi_stmt_1410_req_1 : boolean;
  signal phi_stmt_1410_req_0 : boolean;
  signal phi_stmt_1410_ack_0 : boolean;
  signal ADD_u16_u16_1414_inst_req_0 : boolean;
  signal ADD_u16_u16_1414_inst_ack_0 : boolean;
  signal ADD_u16_u16_1414_inst_req_1 : boolean;
  signal ADD_u16_u16_1414_inst_ack_1 : boolean;
  signal nactive_addr_offset_1439_1415_buf_req_0 : boolean;
  signal nactive_addr_offset_1439_1415_buf_ack_0 : boolean;
  signal nactive_addr_offset_1439_1415_buf_req_1 : boolean;
  signal nactive_addr_offset_1439_1415_buf_ack_1 : boolean;
  signal RPIPE_nic_rx_to_packet_1418_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1418_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1418_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_1418_inst_ack_1 : boolean;
  signal call_stmt_1462_call_req_0 : boolean;
  signal call_stmt_1462_call_ack_0 : boolean;
  signal call_stmt_1462_call_req_1 : boolean;
  signal call_stmt_1462_call_ack_1 : boolean;
  signal do_while_stmt_1408_branch_ack_0 : boolean;
  signal do_while_stmt_1408_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= tag;
  tag_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(23 downto 8) <= max_addr_offset;
  max_addr_offset_buffer <= in_buffer_data_out(23 downto 8);
  in_buffer_data_in(87 downto 24) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(87 downto 24);
  in_buffer_data_in(103 downto 88) <= addr_offset;
  addr_offset_buffer <= in_buffer_data_out(103 downto 88);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_2095_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 20) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(10 downto 0) <= packet_size_11_buffer;
  packet_size_11 <= out_buffer_data_out(10 downto 0);
  out_buffer_data_in(11 downto 11) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(11 downto 11);
  out_buffer_data_in(19 downto 12) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(19 downto 12);
  out_buffer_data_in(tag_length + 19 downto 20) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 19 downto 20);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_2095_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_2095_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_2095_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_2095: Block -- control-path 
    signal writePayloadToMem_CP_2095_elements: BooleanArray(48 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_2095_elements(0) <= writePayloadToMem_CP_2095_start;
    writePayloadToMem_CP_2095_symbol <= writePayloadToMem_CP_2095_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1399/$entry
      -- CP-element group 0: 	 branch_block_stmt_1399/branch_block_stmt_1399__entry__
      -- CP-element group 0: 	 branch_block_stmt_1399/assign_stmt_1407__entry__
      -- CP-element group 0: 	 branch_block_stmt_1399/assign_stmt_1407__exit__
      -- CP-element group 0: 	 branch_block_stmt_1399/do_while_stmt_1408__entry__
      -- CP-element group 0: 	 branch_block_stmt_1399/assign_stmt_1407/$entry
      -- CP-element group 0: 	 branch_block_stmt_1399/assign_stmt_1407/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	48 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1399/$exit
      -- CP-element group 1: 	 branch_block_stmt_1399/branch_block_stmt_1399__exit__
      -- CP-element group 1: 	 branch_block_stmt_1399/do_while_stmt_1408__exit__
      -- CP-element group 1: 	 assign_stmt_1476_to_assign_stmt_1480/$entry
      -- CP-element group 1: 	 assign_stmt_1476_to_assign_stmt_1480/$exit
      -- 
    writePayloadToMem_CP_2095_elements(1) <= writePayloadToMem_CP_2095_elements(48);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1399/do_while_stmt_1408/$entry
      -- CP-element group 2: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408__entry__
      -- 
    writePayloadToMem_CP_2095_elements(2) <= writePayloadToMem_CP_2095_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	48 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408__exit__
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_back
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	47 
    -- CP-element group 5: 	46 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1399/do_while_stmt_1408/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_taken/$entry
      -- 
    writePayloadToMem_CP_2095_elements(5) <= writePayloadToMem_CP_2095_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	45 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_body_done
      -- 
    writePayloadToMem_CP_2095_elements(6) <= writePayloadToMem_CP_2095_elements(45);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/back_edge_to_loop_body
      -- 
    writePayloadToMem_CP_2095_elements(7) <= writePayloadToMem_CP_2095_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/first_time_through_loop_body
      -- 
    writePayloadToMem_CP_2095_elements(8) <= writePayloadToMem_CP_2095_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	44 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1416_sample_start_
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	44 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/condition_evaluated
      -- 
    condition_evaluated_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(10), ack => do_while_stmt_1408_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(15) & writePayloadToMem_CP_2095_elements(44);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	36 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_sample_start__ps
      -- 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(16) & writePayloadToMem_CP_2095_elements(9) & writePayloadToMem_CP_2095_elements(15);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	38 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	45 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1416_sample_completed_
      -- 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(18) & writePayloadToMem_CP_2095_elements(38);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	45 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_2095_elements(12), ack => writePayloadToMem_CP_2095_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	35 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	37 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_update_start__ps
      -- 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(17) & writePayloadToMem_CP_2095_elements(35);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	39 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/aggregated_phi_update_ack
      -- 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(19) & writePayloadToMem_CP_2095_elements(39);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_sample_start_
      -- 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(9) & writePayloadToMem_CP_2095_elements(12);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	42 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_update_start_
      -- 
    writePayloadToMem_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(9) & writePayloadToMem_CP_2095_elements(42);
      gj_writePayloadToMem_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_sample_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	40 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_update_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_loopback_trigger
      -- 
    writePayloadToMem_CP_2095_elements(20) <= writePayloadToMem_CP_2095_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_loopback_sample_req
      -- CP-element group 21: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_loopback_sample_req_ps
      -- 
    phi_stmt_1410_loopback_sample_req_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1410_loopback_sample_req_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(21), ack => phi_stmt_1410_req_1); -- 
    -- Element group writePayloadToMem_CP_2095_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_entry_trigger
      -- 
    writePayloadToMem_CP_2095_elements(22) <= writePayloadToMem_CP_2095_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_entry_sample_req
      -- CP-element group 23: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_entry_sample_req_ps
      -- 
    phi_stmt_1410_entry_sample_req_2143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1410_entry_sample_req_2143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(23), ack => phi_stmt_1410_req_0); -- 
    -- Element group writePayloadToMem_CP_2095_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_phi_mux_ack
      -- CP-element group 24: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1410_phi_mux_ack_ps
      -- 
    phi_stmt_1410_phi_mux_ack_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1410_ack_0, ack => writePayloadToMem_CP_2095_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Sample/rr
      -- 
    rr_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(27), ack => ADD_u16_u16_1414_inst_req_0); -- 
    writePayloadToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(25) & writePayloadToMem_CP_2095_elements(29);
      gj_writePayloadToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Update/cr
      -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(28), ack => ADD_u16_u16_1414_inst_req_1); -- 
    writePayloadToMem_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(26) & writePayloadToMem_CP_2095_elements(30);
      gj_writePayloadToMem_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Sample/ra
      -- 
    ra_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1414_inst_ack_0, ack => writePayloadToMem_CP_2095_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/ADD_u16_u16_1414_Update/ca
      -- 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_1414_inst_ack_1, ack => writePayloadToMem_CP_2095_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Sample/req
      -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(31), ack => nactive_addr_offset_1439_1415_buf_req_0); -- 
    -- Element group writePayloadToMem_CP_2095_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Update/req
      -- 
    req_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(32), ack => nactive_addr_offset_1439_1415_buf_req_1); -- 
    -- Element group writePayloadToMem_CP_2095_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Sample/ack
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nactive_addr_offset_1439_1415_buf_ack_0, ack => writePayloadToMem_CP_2095_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/R_nactive_addr_offset_1415_Update/ack
      -- 
    ack_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nactive_addr_offset_1439_1415_buf_ack_1, ack => writePayloadToMem_CP_2095_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	42 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	14 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1416_update_start_
      -- 
    writePayloadToMem_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(9) & writePayloadToMem_CP_2095_elements(42);
      gj_writePayloadToMem_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	39 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Sample/rr
      -- 
    rr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(36), ack => RPIPE_nic_rx_to_packet_1418_inst_req_0); -- 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(11) & writePayloadToMem_CP_2095_elements(39);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	38 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Update/cr
      -- 
    cr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(37), ack => RPIPE_nic_rx_to_packet_1418_inst_req_1); -- 
    writePayloadToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(14) & writePayloadToMem_CP_2095_elements(38);
      gj_writePayloadToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38: 	37 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Sample/ra
      -- 
    ra_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1418_inst_ack_0, ack => writePayloadToMem_CP_2095_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	15 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	36 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/phi_stmt_1416_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/RPIPE_nic_rx_to_packet_1418_Update/ca
      -- 
    ca_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1418_inst_ack_1, ack => writePayloadToMem_CP_2095_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	19 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Sample/crr
      -- 
    crr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(40), ack => call_stmt_1462_call_req_0); -- 
    writePayloadToMem_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(19) & writePayloadToMem_CP_2095_elements(39);
      gj_writePayloadToMem_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Update/ccr
      -- 
    ccr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_2095_elements(41), ack => call_stmt_1462_call_req_1); -- 
    writePayloadToMem_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_2095_elements(43);
      gj_writePayloadToMem_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	17 
    -- CP-element group 42: 	35 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Sample/cra
      -- 
    cra_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1462_call_ack_0, ack => writePayloadToMem_CP_2095_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/call_stmt_1462_Update/cca
      -- 
    cca_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1462_call_ack_1, ack => writePayloadToMem_CP_2095_elements(43)); -- 
    -- CP-element group 44:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	9 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	10 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writePayloadToMem_CP_2095_elements(44) is a control-delay.
    cp_element_44_delay: control_delay_element  generic map(name => " 44_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_2095_elements(9), ack => writePayloadToMem_CP_2095_elements(44), clk => clk, reset =>reset);
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	12 
    -- CP-element group 45: 	13 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	6 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1399/do_while_stmt_1408/do_while_stmt_1408_loop_body/$exit
      -- 
    writePayloadToMem_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_2095_elements(12) & writePayloadToMem_CP_2095_elements(13) & writePayloadToMem_CP_2095_elements(43);
      gj_writePayloadToMem_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	5 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_exit/$exit
      -- CP-element group 46: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_exit/ack
      -- 
    ack_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1408_branch_ack_0, ack => writePayloadToMem_CP_2095_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	5 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_taken/$exit
      -- CP-element group 47: 	 branch_block_stmt_1399/do_while_stmt_1408/loop_taken/ack
      -- 
    ack_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1408_branch_ack_1, ack => writePayloadToMem_CP_2095_elements(47)); -- 
    -- CP-element group 48:  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	3 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	1 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1399/do_while_stmt_1408/$exit
      -- 
    writePayloadToMem_CP_2095_elements(48) <= writePayloadToMem_CP_2095_elements(3);
    writePayloadToMem_do_while_stmt_1408_terminator_2226: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_1408_terminator_2226", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_2095_elements(6),loop_continue => writePayloadToMem_CP_2095_elements(47),loop_terminate => writePayloadToMem_CP_2095_elements(46),loop_back => writePayloadToMem_CP_2095_elements(4),loop_exit => writePayloadToMem_CP_2095_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1410_phi_seq_2184_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_2095_elements(22);
      writePayloadToMem_CP_2095_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_2095_elements(29);
      writePayloadToMem_CP_2095_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_2095_elements(30);
      writePayloadToMem_CP_2095_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_2095_elements(20);
      writePayloadToMem_CP_2095_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_2095_elements(33);
      writePayloadToMem_CP_2095_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_2095_elements(34);
      writePayloadToMem_CP_2095_elements(21) <= phi_mux_reqs(1);
      phi_stmt_1410_phi_seq_2184 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1410_phi_seq_2184") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_2095_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_2095_elements(18), 
          phi_update_req => writePayloadToMem_CP_2095_elements(14), 
          phi_update_ack => writePayloadToMem_CP_2095_elements(19), 
          phi_mux_ack => writePayloadToMem_CP_2095_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2125_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_2095_elements(7);
        preds(1)  <= writePayloadToMem_CP_2095_elements(8);
        entry_tmerge_2125 : transition_merge -- 
          generic map(name => " entry_tmerge_2125")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_2095_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1414_wire : std_logic_vector(15 downto 0);
    signal AND_u1_u1_1474_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_1445_wire : std_logic_vector(0 downto 0);
    signal EQ_u64_u1_1470_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1473_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1442_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1450_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1452_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_1418_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_1469_wire_constant : std_logic_vector(63 downto 0);
    signal R_WRITEMEM_1456_wire_constant : std_logic_vector(0 downto 0);
    signal SHL_u8_u8_1403_wire : std_logic_vector(7 downto 0);
    signal active_addr_offset_1410 : std_logic_vector(15 downto 0);
    signal continue_flag_1454 : std_logic_vector(0 downto 0);
    signal ignore_return_1462 : std_logic_vector(63 downto 0);
    signal konst_1402_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1413_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1437_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1472_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_1423 : std_logic_vector(0 downto 0);
    signal nactive_addr_offset_1439 : std_logic_vector(15 downto 0);
    signal nactive_addr_offset_1439_1415_buffered : std_logic_vector(15 downto 0);
    signal overflow_1447 : std_logic_vector(0 downto 0);
    signal payloadTag_1407 : std_logic_vector(7 downto 0);
    signal payload_data_1416 : std_logic_vector(72 downto 0);
    signal type_cast_1405_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1459_wire : std_logic_vector(63 downto 0);
    signal wdata_1427 : std_logic_vector(63 downto 0);
    signal wkeep_1431 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_1469_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    R_WRITEMEM_1456_wire_constant <= "0";
    konst_1402_wire_constant <= "00000010";
    konst_1413_wire_constant <= "0000000000001000";
    konst_1437_wire_constant <= "0000000000001000";
    konst_1472_wire_constant <= "00000000";
    type_cast_1405_wire_constant <= "00000010";
    phi_stmt_1410: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u16_u16_1414_wire & nactive_addr_offset_1439_1415_buffered;
      req <= phi_stmt_1410_req_0 & phi_stmt_1410_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1410",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1410_ack_0,
          idata => idata,
          odata => active_addr_offset_1410,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1410
    -- flow-through slice operator slice_1422_inst
    last_bit_1423 <= payload_data_1416(72 downto 72);
    -- flow-through slice operator slice_1426_inst
    wdata_1427 <= payload_data_1416(71 downto 8);
    -- flow-through slice operator slice_1430_inst
    wkeep_1431 <= payload_data_1416(7 downto 0);
    -- interlock W_last_keep_1432_inst
    process(wkeep_1431) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_1431(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    nactive_addr_offset_1439_1415_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nactive_addr_offset_1439_1415_buf_req_0;
      nactive_addr_offset_1439_1415_buf_ack_0<= wack(0);
      rreq(0) <= nactive_addr_offset_1439_1415_buf_req_1;
      nactive_addr_offset_1439_1415_buf_ack_1<= rack(0);
      nactive_addr_offset_1439_1415_buf : InterlockBuffer generic map ( -- 
        name => "nactive_addr_offset_1439_1415_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nactive_addr_offset_1439,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nactive_addr_offset_1439_1415_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1416
    process(RPIPE_nic_rx_to_packet_1418_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_1418_wire(72 downto 0);
      payload_data_1416 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1459_inst
    process(active_addr_offset_1410) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := active_addr_offset_1410(15 downto 0);
      type_cast_1459_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1479_inst
    process(active_addr_offset_1410) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := active_addr_offset_1410(10 downto 0);
      packet_size_11_buffer <= tmp_var; -- 
    end process;
    do_while_stmt_1408_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_1454;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1408_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1408_branch_req_0,
          ack0 => do_while_stmt_1408_branch_ack_0,
          ack1 => do_while_stmt_1408_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u16_u16_1414_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_offset_buffer;
      ADD_u16_u16_1414_wire <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_1414_inst_req_0;
      ADD_u16_u16_1414_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_1414_inst_req_1;
      ADD_u16_u16_1414_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- flow through binary operator ADD_u16_u16_1438_inst
    nactive_addr_offset_1439 <= std_logic_vector(unsigned(active_addr_offset_1410) + unsigned(konst_1437_wire_constant));
    -- flow through binary operator AND_u1_u1_1446_inst
    overflow_1447 <= (NOT_u1_u1_1442_wire and EQ_u16_u1_1445_wire);
    -- flow through binary operator AND_u1_u1_1453_inst
    continue_flag_1454 <= (NOT_u1_u1_1450_wire and NOT_u1_u1_1452_wire);
    -- flow through binary operator AND_u1_u1_1474_inst
    AND_u1_u1_1474_wire <= (EQ_u64_u1_1470_wire and EQ_u8_u1_1473_wire);
    -- flow through binary operator EQ_u16_u1_1445_inst
    process(active_addr_offset_1410, max_addr_offset_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_addr_offset_1410, max_addr_offset_buffer, tmp_var);
      EQ_u16_u1_1445_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u64_u1_1470_inst
    process(wdata_1427) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_1427, R_BAD_PACKET_DATA_1469_wire_constant, tmp_var);
      EQ_u64_u1_1470_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u8_u1_1473_inst
    process(last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_keep_buffer, konst_1472_wire_constant, tmp_var);
      EQ_u8_u1_1473_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1442_inst
    process(last_bit_1423) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_1423, tmp_var);
      NOT_u1_u1_1442_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1450_inst
    process(overflow_1447) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", overflow_1447, tmp_var);
      NOT_u1_u1_1450_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1452_inst
    process(last_bit_1423) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_1423, tmp_var);
      NOT_u1_u1_1452_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_1475_inst
    bad_packet_identifier_buffer <= (overflow_1447 or AND_u1_u1_1474_wire);
    -- flow through binary operator OR_u8_u8_1406_inst
    payloadTag_1407 <= (SHL_u8_u8_1403_wire or type_cast_1405_wire_constant);
    -- flow through binary operator SHL_u8_u8_1403_inst
    process(tag_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tag_buffer, konst_1402_wire_constant, tmp_var);
      SHL_u8_u8_1403_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_1418_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_1418_inst_req_0;
      RPIPE_nic_rx_to_packet_1418_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_1418_inst_req_1;
      RPIPE_nic_rx_to_packet_1418_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_1418_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1462_call 
    accessMemoryDword_call_group_0: Block -- 
      signal data_in: std_logic_vector(200 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 38);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1462_call_req_0;
      call_stmt_1462_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1462_call_req_1;
      call_stmt_1462_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemoryDword_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemoryDword_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= payloadTag_1407 & R_WRITEMEM_1456_wire_constant & base_buf_pointer_buffer & type_cast_1459_wire & wdata_1427;
      ignore_return_1462 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 201,
        owidth => 201,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemoryDword_call_reqs(0),
          ackR => accessMemoryDword_call_acks(0),
          dataR => accessMemoryDword_call_data(200 downto 0),
          tagR => accessMemoryDword_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemoryDword_return_acks(0), -- cross-over
          ackL => accessMemoryDword_return_reqs(0), -- cross-over
          dataL => accessMemoryDword_return_data(63 downto 0),
          tagL => accessMemoryDword_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_lib;
use nic_lib.nic_global_package.all;
entity nic is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    AFB_NIC_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
    AFB_NIC_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MAC_ENABLE: out std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NIC_DEBUG_SIGNAL: out std_logic_vector(255 downto 0);
    NIC_INTR: out std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    RX_ACTIVITY_LOGGER_pipe_read_data: out std_logic_vector(7 downto 0);
    RX_ACTIVITY_LOGGER_pipe_read_req : in std_logic_vector(0 downto 0);
    RX_ACTIVITY_LOGGER_pipe_read_ack : out std_logic_vector(0 downto 0);
    TX_ACTIVITY_LOGGER_pipe_read_data: out std_logic_vector(7 downto 0);
    TX_ACTIVITY_LOGGER_pipe_read_req : in std_logic_vector(0 downto 0);
    TX_ACTIVITY_LOGGER_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data: in std_logic_vector(72 downto 0);
    mac_to_nic_data_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture nic_arch  of nic is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(7 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      S_CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(7 downto 0);
      RX_ACTIVITY_LOGGER_pipe_write_req : out  std_logic_vector(0 downto 0);
      RX_ACTIVITY_LOGGER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      RX_ACTIVITY_LOGGER_pipe_write_data : out  std_logic_vector(7 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(17 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(64 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(87 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(71 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module accessMemoryBase
  component accessMemoryBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      request : in  std_logic_vector(109 downto 0);
      response : out  std_logic_vector(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_DEBUG_SIGNAL_pipe_write_data : out  std_logic_vector(255 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryBase
  signal accessMemoryBase_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryBase_request :  std_logic_vector(109 downto 0);
  signal accessMemoryBase_response :  std_logic_vector(64 downto 0);
  signal accessMemoryBase_in_args    : std_logic_vector(117 downto 0);
  signal accessMemoryBase_out_args   : std_logic_vector(64 downto 0);
  signal accessMemoryBase_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessMemoryBase_tag_out   : std_logic_vector(2 downto 0);
  signal accessMemoryBase_start_req : std_logic;
  signal accessMemoryBase_start_ack : std_logic;
  signal accessMemoryBase_fin_req   : std_logic;
  signal accessMemoryBase_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryBase
  signal accessMemoryBase_call_reqs: std_logic_vector(2 downto 0);
  signal accessMemoryBase_call_acks: std_logic_vector(2 downto 0);
  signal accessMemoryBase_return_reqs: std_logic_vector(2 downto 0);
  signal accessMemoryBase_return_acks: std_logic_vector(2 downto 0);
  signal accessMemoryBase_call_data: std_logic_vector(353 downto 0);
  signal accessMemoryBase_call_tag: std_logic_vector(2 downto 0);
  signal accessMemoryBase_return_data: std_logic_vector(194 downto 0);
  signal accessMemoryBase_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module accessMemoryByte
  component accessMemoryByte is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      byte_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wbyte : in  std_logic_vector(7 downto 0);
      rbyte : out  std_logic_vector(7 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryByte
  signal accessMemoryByte_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryByte_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemoryByte_byte_addr_base :  std_logic_vector(63 downto 0);
  signal accessMemoryByte_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryByte_wbyte :  std_logic_vector(7 downto 0);
  signal accessMemoryByte_rbyte :  std_logic_vector(7 downto 0);
  signal accessMemoryByte_in_args    : std_logic_vector(144 downto 0);
  signal accessMemoryByte_out_args   : std_logic_vector(7 downto 0);
  signal accessMemoryByte_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessMemoryByte_tag_out   : std_logic_vector(1 downto 0);
  signal accessMemoryByte_start_req : std_logic;
  signal accessMemoryByte_start_ack : std_logic;
  signal accessMemoryByte_fin_req   : std_logic;
  signal accessMemoryByte_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryByte
  signal accessMemoryByte_call_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryByte_call_acks: std_logic_vector(0 downto 0);
  signal accessMemoryByte_return_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryByte_return_acks: std_logic_vector(0 downto 0);
  signal accessMemoryByte_call_data: std_logic_vector(144 downto 0);
  signal accessMemoryByte_call_tag: std_logic_vector(0 downto 0);
  signal accessMemoryByte_return_data: std_logic_vector(7 downto 0);
  signal accessMemoryByte_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module accessMemoryByteBase
  component accessMemoryByteBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      byte_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wbyte : in  std_logic_vector(7 downto 0);
      rbyte : out  std_logic_vector(7 downto 0);
      calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
      calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
      calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
      calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
      accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
      accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryByteBase
  signal accessMemoryByteBase_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryByteBase_lock :  std_logic_vector(0 downto 0);
  signal accessMemoryByteBase_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemoryByteBase_byte_addr_base :  std_logic_vector(63 downto 0);
  signal accessMemoryByteBase_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryByteBase_wbyte :  std_logic_vector(7 downto 0);
  signal accessMemoryByteBase_rbyte :  std_logic_vector(7 downto 0);
  signal accessMemoryByteBase_in_args    : std_logic_vector(145 downto 0);
  signal accessMemoryByteBase_out_args   : std_logic_vector(7 downto 0);
  signal accessMemoryByteBase_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessMemoryByteBase_tag_out   : std_logic_vector(2 downto 0);
  signal accessMemoryByteBase_start_req : std_logic;
  signal accessMemoryByteBase_start_ack : std_logic;
  signal accessMemoryByteBase_fin_req   : std_logic;
  signal accessMemoryByteBase_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryByteBase
  signal accessMemoryByteBase_call_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryByteBase_call_acks: std_logic_vector(0 downto 0);
  signal accessMemoryByteBase_return_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryByteBase_return_acks: std_logic_vector(0 downto 0);
  signal accessMemoryByteBase_call_data: std_logic_vector(145 downto 0);
  signal accessMemoryByteBase_call_tag: std_logic_vector(1 downto 0);
  signal accessMemoryByteBase_return_data: std_logic_vector(7 downto 0);
  signal accessMemoryByteBase_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemoryDword
  component accessMemoryDword is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryDword
  signal accessMemoryDword_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryDword_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemoryDword_base_addr :  std_logic_vector(63 downto 0);
  signal accessMemoryDword_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryDword_wdata :  std_logic_vector(63 downto 0);
  signal accessMemoryDword_rdata :  std_logic_vector(63 downto 0);
  signal accessMemoryDword_in_args    : std_logic_vector(200 downto 0);
  signal accessMemoryDword_out_args   : std_logic_vector(63 downto 0);
  signal accessMemoryDword_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal accessMemoryDword_tag_out   : std_logic_vector(4 downto 0);
  signal accessMemoryDword_start_req : std_logic;
  signal accessMemoryDword_start_ack : std_logic;
  signal accessMemoryDword_fin_req   : std_logic;
  signal accessMemoryDword_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryDword
  signal accessMemoryDword_call_reqs: std_logic_vector(6 downto 0);
  signal accessMemoryDword_call_acks: std_logic_vector(6 downto 0);
  signal accessMemoryDword_return_reqs: std_logic_vector(6 downto 0);
  signal accessMemoryDword_return_acks: std_logic_vector(6 downto 0);
  signal accessMemoryDword_call_data: std_logic_vector(1406 downto 0);
  signal accessMemoryDword_call_tag: std_logic_vector(13 downto 0);
  signal accessMemoryDword_return_data: std_logic_vector(447 downto 0);
  signal accessMemoryDword_return_tag: std_logic_vector(13 downto 0);
  -- declarations related to module accessMemoryDwordBase
  component accessMemoryDwordBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
      calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
      calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
      calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
      accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
      accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryDwordBase
  signal accessMemoryDwordBase_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryDwordBase_lock :  std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_base_addr :  std_logic_vector(63 downto 0);
  signal accessMemoryDwordBase_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryDwordBase_wdata :  std_logic_vector(63 downto 0);
  signal accessMemoryDwordBase_rdata :  std_logic_vector(63 downto 0);
  signal accessMemoryDwordBase_in_args    : std_logic_vector(201 downto 0);
  signal accessMemoryDwordBase_out_args   : std_logic_vector(63 downto 0);
  signal accessMemoryDwordBase_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessMemoryDwordBase_tag_out   : std_logic_vector(1 downto 0);
  signal accessMemoryDwordBase_start_req : std_logic;
  signal accessMemoryDwordBase_start_ack : std_logic;
  signal accessMemoryDwordBase_fin_req   : std_logic;
  signal accessMemoryDwordBase_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryDwordBase
  signal accessMemoryDwordBase_call_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_call_acks: std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_return_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_return_acks: std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_call_data: std_logic_vector(201 downto 0);
  signal accessMemoryDwordBase_call_tag: std_logic_vector(0 downto 0);
  signal accessMemoryDwordBase_return_data: std_logic_vector(63 downto 0);
  signal accessMemoryDwordBase_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module accessMemoryLdStub
  component accessMemoryLdStub is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      byte_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      rbyte : out  std_logic_vector(7 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryLdStub
  signal accessMemoryLdStub_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryLdStub_byte_addr_base :  std_logic_vector(63 downto 0);
  signal accessMemoryLdStub_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryLdStub_rbyte :  std_logic_vector(7 downto 0);
  signal accessMemoryLdStub_in_args    : std_logic_vector(135 downto 0);
  signal accessMemoryLdStub_out_args   : std_logic_vector(7 downto 0);
  signal accessMemoryLdStub_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessMemoryLdStub_tag_out   : std_logic_vector(1 downto 0);
  signal accessMemoryLdStub_start_req : std_logic;
  signal accessMemoryLdStub_start_ack : std_logic;
  signal accessMemoryLdStub_fin_req   : std_logic;
  signal accessMemoryLdStub_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryLdStub
  signal accessMemoryLdStub_call_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryLdStub_call_acks: std_logic_vector(0 downto 0);
  signal accessMemoryLdStub_return_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryLdStub_return_acks: std_logic_vector(0 downto 0);
  signal accessMemoryLdStub_call_data: std_logic_vector(135 downto 0);
  signal accessMemoryLdStub_call_tag: std_logic_vector(0 downto 0);
  signal accessMemoryLdStub_return_data: std_logic_vector(7 downto 0);
  signal accessMemoryLdStub_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module accessMemoryWord
  component accessMemoryWord is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      doMemAccess_call_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_call_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_call_data : out  std_logic_vector(202 downto 0);
      doMemAccess_call_tag  :  out  std_logic_vector(0 downto 0);
      doMemAccess_return_reqs : out  std_logic_vector(0 downto 0);
      doMemAccess_return_acks : in   std_logic_vector(0 downto 0);
      doMemAccess_return_data : in   std_logic_vector(63 downto 0);
      doMemAccess_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryWord
  signal accessMemoryWord_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryWord_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemoryWord_word_addr_base :  std_logic_vector(63 downto 0);
  signal accessMemoryWord_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryWord_wword :  std_logic_vector(31 downto 0);
  signal accessMemoryWord_rword :  std_logic_vector(31 downto 0);
  signal accessMemoryWord_in_args    : std_logic_vector(168 downto 0);
  signal accessMemoryWord_out_args   : std_logic_vector(31 downto 0);
  signal accessMemoryWord_tag_in    : std_logic_vector(3 downto 0) := (others => '0');
  signal accessMemoryWord_tag_out   : std_logic_vector(3 downto 0);
  signal accessMemoryWord_start_req : std_logic;
  signal accessMemoryWord_start_ack : std_logic;
  signal accessMemoryWord_fin_req   : std_logic;
  signal accessMemoryWord_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryWord
  signal accessMemoryWord_call_reqs: std_logic_vector(5 downto 0);
  signal accessMemoryWord_call_acks: std_logic_vector(5 downto 0);
  signal accessMemoryWord_return_reqs: std_logic_vector(5 downto 0);
  signal accessMemoryWord_return_acks: std_logic_vector(5 downto 0);
  signal accessMemoryWord_call_data: std_logic_vector(1013 downto 0);
  signal accessMemoryWord_call_tag: std_logic_vector(5 downto 0);
  signal accessMemoryWord_return_data: std_logic_vector(191 downto 0);
  signal accessMemoryWord_return_tag: std_logic_vector(5 downto 0);
  -- declarations related to module accessMemoryWordBase
  component accessMemoryWordBase is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      word_addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wword : in  std_logic_vector(31 downto 0);
      rword : out  std_logic_vector(31 downto 0);
      calculateAddress36_call_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_call_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_call_data : out  std_logic_vector(127 downto 0);
      calculateAddress36_call_tag  :  out  std_logic_vector(0 downto 0);
      calculateAddress36_return_reqs : out  std_logic_vector(0 downto 0);
      calculateAddress36_return_acks : in   std_logic_vector(0 downto 0);
      calculateAddress36_return_data : in   std_logic_vector(35 downto 0);
      calculateAddress36_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_call_data : out  std_logic_vector(117 downto 0);
      accessMemoryBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryBase_return_data : in   std_logic_vector(64 downto 0);
      accessMemoryBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemoryWordBase
  signal accessMemoryWordBase_tag :  std_logic_vector(7 downto 0);
  signal accessMemoryWordBase_lock :  std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_word_addr_base :  std_logic_vector(63 downto 0);
  signal accessMemoryWordBase_offset :  std_logic_vector(63 downto 0);
  signal accessMemoryWordBase_wword :  std_logic_vector(31 downto 0);
  signal accessMemoryWordBase_rword :  std_logic_vector(31 downto 0);
  signal accessMemoryWordBase_in_args    : std_logic_vector(169 downto 0);
  signal accessMemoryWordBase_out_args   : std_logic_vector(31 downto 0);
  signal accessMemoryWordBase_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessMemoryWordBase_tag_out   : std_logic_vector(1 downto 0);
  signal accessMemoryWordBase_start_req : std_logic;
  signal accessMemoryWordBase_start_ack : std_logic;
  signal accessMemoryWordBase_fin_req   : std_logic;
  signal accessMemoryWordBase_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemoryWordBase
  signal accessMemoryWordBase_call_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_call_acks: std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_return_reqs: std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_return_acks: std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_call_data: std_logic_vector(169 downto 0);
  signal accessMemoryWordBase_call_tag: std_logic_vector(0 downto 0);
  signal accessMemoryWordBase_return_data: std_logic_vector(31 downto 0);
  signal accessMemoryWordBase_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module accessQueueElement
  component accessQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      index : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessQueueElement
  signal accessQueueElement_tag :  std_logic_vector(7 downto 0);
  signal accessQueueElement_rwbar :  std_logic_vector(0 downto 0);
  signal accessQueueElement_base_addr :  std_logic_vector(63 downto 0);
  signal accessQueueElement_index :  std_logic_vector(31 downto 0);
  signal accessQueueElement_wdata :  std_logic_vector(63 downto 0);
  signal accessQueueElement_rdata :  std_logic_vector(63 downto 0);
  signal accessQueueElement_in_args    : std_logic_vector(168 downto 0);
  signal accessQueueElement_out_args   : std_logic_vector(63 downto 0);
  signal accessQueueElement_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessQueueElement_tag_out   : std_logic_vector(2 downto 0);
  signal accessQueueElement_start_req : std_logic;
  signal accessQueueElement_start_ack : std_logic;
  signal accessQueueElement_fin_req   : std_logic;
  signal accessQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module accessQueueElement
  signal accessQueueElement_call_reqs: std_logic_vector(1 downto 0);
  signal accessQueueElement_call_acks: std_logic_vector(1 downto 0);
  signal accessQueueElement_return_reqs: std_logic_vector(1 downto 0);
  signal accessQueueElement_return_acks: std_logic_vector(1 downto 0);
  signal accessQueueElement_call_data: std_logic_vector(337 downto 0);
  signal accessQueueElement_call_tag: std_logic_vector(1 downto 0);
  signal accessQueueElement_return_data: std_logic_vector(127 downto 0);
  signal accessQueueElement_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessQueueLength
  component accessQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessQueueLength
  signal accessQueueLength_tag :  std_logic_vector(7 downto 0);
  signal accessQueueLength_rwbar :  std_logic_vector(0 downto 0);
  signal accessQueueLength_qptr :  std_logic_vector(63 downto 0);
  signal accessQueueLength_wdata :  std_logic_vector(31 downto 0);
  signal accessQueueLength_rdata :  std_logic_vector(31 downto 0);
  signal accessQueueLength_in_args    : std_logic_vector(104 downto 0);
  signal accessQueueLength_out_args   : std_logic_vector(31 downto 0);
  signal accessQueueLength_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessQueueLength_tag_out   : std_logic_vector(1 downto 0);
  signal accessQueueLength_start_req : std_logic;
  signal accessQueueLength_start_ack : std_logic;
  signal accessQueueLength_fin_req   : std_logic;
  signal accessQueueLength_fin_ack : std_logic;
  -- caller side aggregated signals for module accessQueueLength
  signal accessQueueLength_call_reqs: std_logic_vector(0 downto 0);
  signal accessQueueLength_call_acks: std_logic_vector(0 downto 0);
  signal accessQueueLength_return_reqs: std_logic_vector(0 downto 0);
  signal accessQueueLength_return_acks: std_logic_vector(0 downto 0);
  signal accessQueueLength_call_data: std_logic_vector(104 downto 0);
  signal accessQueueLength_call_tag: std_logic_vector(0 downto 0);
  signal accessQueueLength_return_data: std_logic_vector(31 downto 0);
  signal accessQueueLength_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module accessQueueMisc
  component accessQueueMisc is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessQueueMisc
  signal accessQueueMisc_tag :  std_logic_vector(7 downto 0);
  signal accessQueueMisc_rwbar :  std_logic_vector(0 downto 0);
  signal accessQueueMisc_qptr :  std_logic_vector(63 downto 0);
  signal accessQueueMisc_wdata :  std_logic_vector(31 downto 0);
  signal accessQueueMisc_rdata :  std_logic_vector(31 downto 0);
  signal accessQueueMisc_in_args    : std_logic_vector(104 downto 0);
  signal accessQueueMisc_out_args   : std_logic_vector(31 downto 0);
  signal accessQueueMisc_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessQueueMisc_tag_out   : std_logic_vector(1 downto 0);
  signal accessQueueMisc_start_req : std_logic;
  signal accessQueueMisc_start_ack : std_logic;
  signal accessQueueMisc_fin_req   : std_logic;
  signal accessQueueMisc_fin_ack : std_logic;
  -- caller side aggregated signals for module accessQueueMisc
  signal accessQueueMisc_call_reqs: std_logic_vector(0 downto 0);
  signal accessQueueMisc_call_acks: std_logic_vector(0 downto 0);
  signal accessQueueMisc_return_reqs: std_logic_vector(0 downto 0);
  signal accessQueueMisc_return_acks: std_logic_vector(0 downto 0);
  signal accessQueueMisc_call_data: std_logic_vector(104 downto 0);
  signal accessQueueMisc_call_tag: std_logic_vector(0 downto 0);
  signal accessQueueMisc_return_data: std_logic_vector(31 downto 0);
  signal accessQueueMisc_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module accessQueueReadIndex
  component accessQueueReadIndex is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessQueueReadIndex
  signal accessQueueReadIndex_tag :  std_logic_vector(7 downto 0);
  signal accessQueueReadIndex_rwbar :  std_logic_vector(0 downto 0);
  signal accessQueueReadIndex_qptr :  std_logic_vector(63 downto 0);
  signal accessQueueReadIndex_wdata :  std_logic_vector(31 downto 0);
  signal accessQueueReadIndex_rdata :  std_logic_vector(31 downto 0);
  signal accessQueueReadIndex_in_args    : std_logic_vector(104 downto 0);
  signal accessQueueReadIndex_out_args   : std_logic_vector(31 downto 0);
  signal accessQueueReadIndex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessQueueReadIndex_tag_out   : std_logic_vector(2 downto 0);
  signal accessQueueReadIndex_start_req : std_logic;
  signal accessQueueReadIndex_start_ack : std_logic;
  signal accessQueueReadIndex_fin_req   : std_logic;
  signal accessQueueReadIndex_fin_ack : std_logic;
  -- caller side aggregated signals for module accessQueueReadIndex
  signal accessQueueReadIndex_call_reqs: std_logic_vector(1 downto 0);
  signal accessQueueReadIndex_call_acks: std_logic_vector(1 downto 0);
  signal accessQueueReadIndex_return_reqs: std_logic_vector(1 downto 0);
  signal accessQueueReadIndex_return_acks: std_logic_vector(1 downto 0);
  signal accessQueueReadIndex_call_data: std_logic_vector(209 downto 0);
  signal accessQueueReadIndex_call_tag: std_logic_vector(1 downto 0);
  signal accessQueueReadIndex_return_data: std_logic_vector(63 downto 0);
  signal accessQueueReadIndex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessQueueTotalMsgs
  component accessQueueTotalMsgs is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessQueueTotalMsgs
  signal accessQueueTotalMsgs_tag :  std_logic_vector(7 downto 0);
  signal accessQueueTotalMsgs_rwbar :  std_logic_vector(0 downto 0);
  signal accessQueueTotalMsgs_qptr :  std_logic_vector(63 downto 0);
  signal accessQueueTotalMsgs_wdata :  std_logic_vector(31 downto 0);
  signal accessQueueTotalMsgs_rdata :  std_logic_vector(31 downto 0);
  signal accessQueueTotalMsgs_in_args    : std_logic_vector(104 downto 0);
  signal accessQueueTotalMsgs_out_args   : std_logic_vector(31 downto 0);
  signal accessQueueTotalMsgs_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessQueueTotalMsgs_tag_out   : std_logic_vector(2 downto 0);
  signal accessQueueTotalMsgs_start_req : std_logic;
  signal accessQueueTotalMsgs_start_ack : std_logic;
  signal accessQueueTotalMsgs_fin_req   : std_logic;
  signal accessQueueTotalMsgs_fin_ack : std_logic;
  -- caller side aggregated signals for module accessQueueTotalMsgs
  signal accessQueueTotalMsgs_call_reqs: std_logic_vector(1 downto 0);
  signal accessQueueTotalMsgs_call_acks: std_logic_vector(1 downto 0);
  signal accessQueueTotalMsgs_return_reqs: std_logic_vector(1 downto 0);
  signal accessQueueTotalMsgs_return_acks: std_logic_vector(1 downto 0);
  signal accessQueueTotalMsgs_call_data: std_logic_vector(209 downto 0);
  signal accessQueueTotalMsgs_call_tag: std_logic_vector(1 downto 0);
  signal accessQueueTotalMsgs_return_data: std_logic_vector(63 downto 0);
  signal accessQueueTotalMsgs_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessQueueWriteIndex
  component accessQueueWriteIndex is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      qptr : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessQueueWriteIndex
  signal accessQueueWriteIndex_tag :  std_logic_vector(7 downto 0);
  signal accessQueueWriteIndex_rwbar :  std_logic_vector(0 downto 0);
  signal accessQueueWriteIndex_qptr :  std_logic_vector(63 downto 0);
  signal accessQueueWriteIndex_wdata :  std_logic_vector(31 downto 0);
  signal accessQueueWriteIndex_rdata :  std_logic_vector(31 downto 0);
  signal accessQueueWriteIndex_in_args    : std_logic_vector(104 downto 0);
  signal accessQueueWriteIndex_out_args   : std_logic_vector(31 downto 0);
  signal accessQueueWriteIndex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessQueueWriteIndex_tag_out   : std_logic_vector(2 downto 0);
  signal accessQueueWriteIndex_start_req : std_logic;
  signal accessQueueWriteIndex_start_ack : std_logic;
  signal accessQueueWriteIndex_fin_req   : std_logic;
  signal accessQueueWriteIndex_fin_ack : std_logic;
  -- caller side aggregated signals for module accessQueueWriteIndex
  signal accessQueueWriteIndex_call_reqs: std_logic_vector(1 downto 0);
  signal accessQueueWriteIndex_call_acks: std_logic_vector(1 downto 0);
  signal accessQueueWriteIndex_return_reqs: std_logic_vector(1 downto 0);
  signal accessQueueWriteIndex_return_acks: std_logic_vector(1 downto 0);
  signal accessQueueWriteIndex_call_data: std_logic_vector(209 downto 0);
  signal accessQueueWriteIndex_call_tag: std_logic_vector(1 downto 0);
  signal accessQueueWriteIndex_return_data: std_logic_vector(63 downto 0);
  signal accessQueueWriteIndex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessRegister
  component accessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      index : in  std_logic_vector(7 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessRegister
  signal accessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal accessRegister_bmask :  std_logic_vector(3 downto 0);
  signal accessRegister_index :  std_logic_vector(7 downto 0);
  signal accessRegister_wdata :  std_logic_vector(31 downto 0);
  signal accessRegister_rdata :  std_logic_vector(31 downto 0);
  signal accessRegister_in_args    : std_logic_vector(44 downto 0);
  signal accessRegister_out_args   : std_logic_vector(31 downto 0);
  signal accessRegister_tag_in    : std_logic_vector(5 downto 0) := (others => '0');
  signal accessRegister_tag_out   : std_logic_vector(5 downto 0);
  signal accessRegister_start_req : std_logic;
  signal accessRegister_start_ack : std_logic;
  signal accessRegister_fin_req   : std_logic;
  signal accessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module accessRegister
  signal accessRegister_call_reqs: std_logic_vector(9 downto 0);
  signal accessRegister_call_acks: std_logic_vector(9 downto 0);
  signal accessRegister_return_reqs: std_logic_vector(9 downto 0);
  signal accessRegister_return_acks: std_logic_vector(9 downto 0);
  signal accessRegister_call_data: std_logic_vector(449 downto 0);
  signal accessRegister_call_tag: std_logic_vector(19 downto 0);
  signal accessRegister_return_data: std_logic_vector(319 downto 0);
  signal accessRegister_return_tag: std_logic_vector(19 downto 0);
  -- declarations related to module acquireLock
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock_address_pointer : in  std_logic_vector(63 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryLdStub_call_data : out  std_logic_vector(135 downto 0);
      accessMemoryLdStub_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryLdStub_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryLdStub_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireLock
  signal acquireLock_tag :  std_logic_vector(7 downto 0);
  signal acquireLock_lock_address_pointer :  std_logic_vector(63 downto 0);
  signal acquireLock_m_ok :  std_logic_vector(0 downto 0);
  signal acquireLock_in_args    : std_logic_vector(71 downto 0);
  signal acquireLock_out_args   : std_logic_vector(0 downto 0);
  signal acquireLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireLock_tag_out   : std_logic_vector(2 downto 0);
  signal acquireLock_start_req : std_logic;
  signal acquireLock_start_ack : std_logic;
  signal acquireLock_fin_req   : std_logic;
  signal acquireLock_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireLock
  signal acquireLock_call_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_call_acks: std_logic_vector(1 downto 0);
  signal acquireLock_return_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_return_acks: std_logic_vector(1 downto 0);
  signal acquireLock_call_data: std_logic_vector(143 downto 0);
  signal acquireLock_call_tag: std_logic_vector(1 downto 0);
  signal acquireLock_return_data: std_logic_vector(1 downto 0);
  signal acquireLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module calculateAddress36
  component calculateAddress36 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr_base : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      addr : out  std_logic_vector(35 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module calculateAddress36
  signal calculateAddress36_addr_base :  std_logic_vector(63 downto 0);
  signal calculateAddress36_offset :  std_logic_vector(63 downto 0);
  signal calculateAddress36_addr :  std_logic_vector(35 downto 0);
  signal calculateAddress36_in_args    : std_logic_vector(127 downto 0);
  signal calculateAddress36_out_args   : std_logic_vector(35 downto 0);
  signal calculateAddress36_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal calculateAddress36_tag_out   : std_logic_vector(2 downto 0);
  signal calculateAddress36_start_req : std_logic;
  signal calculateAddress36_start_ack : std_logic;
  signal calculateAddress36_fin_req   : std_logic;
  signal calculateAddress36_fin_ack : std_logic;
  -- caller side aggregated signals for module calculateAddress36
  signal calculateAddress36_call_reqs: std_logic_vector(2 downto 0);
  signal calculateAddress36_call_acks: std_logic_vector(2 downto 0);
  signal calculateAddress36_return_reqs: std_logic_vector(2 downto 0);
  signal calculateAddress36_return_acks: std_logic_vector(2 downto 0);
  signal calculateAddress36_call_data: std_logic_vector(383 downto 0);
  signal calculateAddress36_call_tag: std_logic_vector(2 downto 0);
  signal calculateAddress36_return_data: std_logic_vector(107 downto 0);
  signal calculateAddress36_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module controlDaemon
  component controlDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      QUEUE_MONITOR_SIGNAL : in std_logic_vector(31 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      NIC_INTR_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_data : out  std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      NIC_INTR_INTERNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_INTERNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_INTERNAL_pipe_write_data : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(1 downto 0);
      accessRegister_call_acks : in   std_logic_vector(1 downto 0);
      accessRegister_call_data : out  std_logic_vector(89 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(1 downto 0);
      accessRegister_return_acks : in   std_logic_vector(1 downto 0);
      accessRegister_return_data : in   std_logic_vector(63 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(3 downto 0);
      setGlobalSignals_call_reqs : out  std_logic_vector(0 downto 0);
      setGlobalSignals_call_acks : in   std_logic_vector(0 downto 0);
      setGlobalSignals_call_tag  :  out  std_logic_vector(0 downto 0);
      setGlobalSignals_return_reqs : out  std_logic_vector(0 downto 0);
      setGlobalSignals_return_acks : in   std_logic_vector(0 downto 0);
      setGlobalSignals_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module controlDaemon
  signal controlDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal controlDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal controlDaemon_start_req : std_logic;
  signal controlDaemon_start_ack : std_logic;
  signal controlDaemon_fin_req   : std_logic;
  signal controlDaemon_fin_ack : std_logic;
  -- declarations related to module delay_time
  -- declarations related to module doMemAccess
  component doMemAccess is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      opcode : in  std_logic_vector(2 downto 0);
      base_addr : in  std_logic_vector(63 downto 0);
      offset : in  std_logic_vector(63 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      memory_access_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      memory_access_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_call_data : out  std_logic_vector(169 downto 0);
      accessMemoryWordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWordBase_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWordBase_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_call_data : out  std_logic_vector(145 downto 0);
      accessMemoryByteBase_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryByteBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByteBase_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByteBase_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemoryDwordBase_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_call_data : out  std_logic_vector(201 downto 0);
      accessMemoryDwordBase_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDwordBase_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDwordBase_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module doMemAccess
  signal doMemAccess_tag :  std_logic_vector(7 downto 0);
  signal doMemAccess_opcode :  std_logic_vector(2 downto 0);
  signal doMemAccess_base_addr :  std_logic_vector(63 downto 0);
  signal doMemAccess_offset :  std_logic_vector(63 downto 0);
  signal doMemAccess_wdata :  std_logic_vector(63 downto 0);
  signal doMemAccess_rdata :  std_logic_vector(63 downto 0);
  signal doMemAccess_in_args    : std_logic_vector(202 downto 0);
  signal doMemAccess_out_args   : std_logic_vector(63 downto 0);
  signal doMemAccess_tag_in    : std_logic_vector(3 downto 0) := (others => '0');
  signal doMemAccess_tag_out   : std_logic_vector(3 downto 0);
  signal doMemAccess_start_req : std_logic;
  signal doMemAccess_start_ack : std_logic;
  signal doMemAccess_fin_req   : std_logic;
  signal doMemAccess_fin_ack : std_logic;
  -- caller side aggregated signals for module doMemAccess
  signal doMemAccess_call_reqs: std_logic_vector(3 downto 0);
  signal doMemAccess_call_acks: std_logic_vector(3 downto 0);
  signal doMemAccess_return_reqs: std_logic_vector(3 downto 0);
  signal doMemAccess_return_acks: std_logic_vector(3 downto 0);
  signal doMemAccess_call_data: std_logic_vector(811 downto 0);
  signal doMemAccess_call_tag: std_logic_vector(3 downto 0);
  signal doMemAccess_return_data: std_logic_vector(255 downto 0);
  signal doMemAccess_return_tag: std_logic_vector(3 downto 0);
  -- declarations related to module getBaseIndex
  -- declarations related to module getQueueBufPointer
  component getQueueBufPointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueBufPointer
  signal getQueueBufPointer_queue_type :  std_logic_vector(1 downto 0);
  signal getQueueBufPointer_server_id :  std_logic_vector(7 downto 0);
  signal getQueueBufPointer_qptr :  std_logic_vector(63 downto 0);
  signal getQueueBufPointer_in_args    : std_logic_vector(9 downto 0);
  signal getQueueBufPointer_out_args   : std_logic_vector(63 downto 0);
  signal getQueueBufPointer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueueBufPointer_tag_out   : std_logic_vector(2 downto 0);
  signal getQueueBufPointer_start_req : std_logic;
  signal getQueueBufPointer_start_ack : std_logic;
  signal getQueueBufPointer_fin_req   : std_logic;
  signal getQueueBufPointer_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueBufPointer
  signal getQueueBufPointer_call_reqs: std_logic_vector(1 downto 0);
  signal getQueueBufPointer_call_acks: std_logic_vector(1 downto 0);
  signal getQueueBufPointer_return_reqs: std_logic_vector(1 downto 0);
  signal getQueueBufPointer_return_acks: std_logic_vector(1 downto 0);
  signal getQueueBufPointer_call_data: std_logic_vector(19 downto 0);
  signal getQueueBufPointer_call_tag: std_logic_vector(1 downto 0);
  signal getQueueBufPointer_return_data: std_logic_vector(127 downto 0);
  signal getQueueBufPointer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      buf_base_addr : in  std_logic_vector(63 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(63 downto 0);
      accessQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_call_data : out  std_logic_vector(168 downto 0);
      accessQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_return_data : in   std_logic_vector(63 downto 0);
      accessQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_tag :  std_logic_vector(7 downto 0);
  signal getQueueElement_buf_base_addr :  std_logic_vector(63 downto 0);
  signal getQueueElement_read_index :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(63 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(103 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(63 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(103 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(63 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueueLength
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      queue_length : out  std_logic_vector(31 downto 0);
      accessQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueLength_call_data : out  std_logic_vector(104 downto 0);
      accessQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueLength_return_data : in   std_logic_vector(31 downto 0);
      accessQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueLength
  signal getQueueLength_tag :  std_logic_vector(7 downto 0);
  signal getQueueLength_q_base_address :  std_logic_vector(63 downto 0);
  signal getQueueLength_queue_length :  std_logic_vector(31 downto 0);
  signal getQueueLength_in_args    : std_logic_vector(71 downto 0);
  signal getQueueLength_out_args   : std_logic_vector(31 downto 0);
  signal getQueueLength_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueueLength_tag_out   : std_logic_vector(2 downto 0);
  signal getQueueLength_start_req : std_logic;
  signal getQueueLength_start_ack : std_logic;
  signal getQueueLength_fin_req   : std_logic;
  signal getQueueLength_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueLength
  signal getQueueLength_call_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_call_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_return_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_return_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_call_data: std_logic_vector(143 downto 0);
  signal getQueueLength_call_tag: std_logic_vector(1 downto 0);
  signal getQueueLength_return_data: std_logic_vector(63 downto 0);
  signal getQueueLength_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueueLockPointer
  component getQueueLockPointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueLockPointer
  signal getQueueLockPointer_queue_type :  std_logic_vector(1 downto 0);
  signal getQueueLockPointer_server_id :  std_logic_vector(7 downto 0);
  signal getQueueLockPointer_qptr :  std_logic_vector(63 downto 0);
  signal getQueueLockPointer_in_args    : std_logic_vector(9 downto 0);
  signal getQueueLockPointer_out_args   : std_logic_vector(63 downto 0);
  signal getQueueLockPointer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueueLockPointer_tag_out   : std_logic_vector(2 downto 0);
  signal getQueueLockPointer_start_req : std_logic;
  signal getQueueLockPointer_start_ack : std_logic;
  signal getQueueLockPointer_fin_req   : std_logic;
  signal getQueueLockPointer_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueLockPointer
  signal getQueueLockPointer_call_reqs: std_logic_vector(1 downto 0);
  signal getQueueLockPointer_call_acks: std_logic_vector(1 downto 0);
  signal getQueueLockPointer_return_reqs: std_logic_vector(1 downto 0);
  signal getQueueLockPointer_return_acks: std_logic_vector(1 downto 0);
  signal getQueueLockPointer_call_data: std_logic_vector(19 downto 0);
  signal getQueueLockPointer_call_tag: std_logic_vector(1 downto 0);
  signal getQueueLockPointer_return_data: std_logic_vector(127 downto 0);
  signal getQueueLockPointer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueuePointer
  component getQueuePointer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      qptr : out  std_logic_vector(63 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointer
  signal getQueuePointer_queue_type :  std_logic_vector(1 downto 0);
  signal getQueuePointer_server_id :  std_logic_vector(7 downto 0);
  signal getQueuePointer_qptr :  std_logic_vector(63 downto 0);
  signal getQueuePointer_in_args    : std_logic_vector(9 downto 0);
  signal getQueuePointer_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointer_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointer_start_req : std_logic;
  signal getQueuePointer_start_ack : std_logic;
  signal getQueuePointer_fin_req   : std_logic;
  signal getQueuePointer_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointer
  signal getQueuePointer_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointer_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointer_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointer_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointer_call_data: std_logic_vector(19 downto 0);
  signal getQueuePointer_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointer_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_tag :  std_logic_vector(7 downto 0);
  signal getQueuePointers_q_base_address :  std_logic_vector(63 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(71 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(143 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTotalMessages
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
      accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTotalMessages
  signal getTotalMessages_tag :  std_logic_vector(7 downto 0);
  signal getTotalMessages_q_base_address :  std_logic_vector(63 downto 0);
  signal getTotalMessages_total_msgs :  std_logic_vector(31 downto 0);
  signal getTotalMessages_in_args    : std_logic_vector(71 downto 0);
  signal getTotalMessages_out_args   : std_logic_vector(31 downto 0);
  signal getTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal getTotalMessages_start_req : std_logic;
  signal getTotalMessages_start_ack : std_logic;
  signal getTotalMessages_fin_req   : std_logic;
  signal getTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module getTotalMessages
  signal getTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_data: std_logic_vector(143 downto 0);
  signal getTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_data: std_logic_vector(63 downto 0);
  signal getTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      server_index : in  std_logic_vector(7 downto 0);
      pkt_pointer : out  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(17 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(64 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_tag :  std_logic_vector(7 downto 0);
  signal getTxPacketPointerFromServer_server_index :  std_logic_vector(7 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(63 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(15 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(64 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(15 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(64 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module incrementNumberOfPacketsReceived
  component incrementNumberOfPacketsReceived is -- 
    generic (tag_length : integer); 
    port ( -- 
      incrementRegister_call_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_call_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_call_data : out  std_logic_vector(7 downto 0);
      incrementRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementRegister_return_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_return_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_return_data : in   std_logic_vector(31 downto 0);
      incrementRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module incrementNumberOfPacketsReceived
  signal incrementNumberOfPacketsReceived_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal incrementNumberOfPacketsReceived_tag_out   : std_logic_vector(1 downto 0);
  signal incrementNumberOfPacketsReceived_start_req : std_logic;
  signal incrementNumberOfPacketsReceived_start_ack : std_logic;
  signal incrementNumberOfPacketsReceived_fin_req   : std_logic;
  signal incrementNumberOfPacketsReceived_fin_ack : std_logic;
  -- caller side aggregated signals for module incrementNumberOfPacketsReceived
  signal incrementNumberOfPacketsReceived_call_reqs: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsReceived_call_acks: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsReceived_return_reqs: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsReceived_return_acks: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsReceived_call_tag: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsReceived_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module incrementNumberOfPacketsTransmitted
  component incrementNumberOfPacketsTransmitted is -- 
    generic (tag_length : integer); 
    port ( -- 
      incrementRegister_call_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_call_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_call_data : out  std_logic_vector(7 downto 0);
      incrementRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementRegister_return_reqs : out  std_logic_vector(0 downto 0);
      incrementRegister_return_acks : in   std_logic_vector(0 downto 0);
      incrementRegister_return_data : in   std_logic_vector(31 downto 0);
      incrementRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module incrementNumberOfPacketsTransmitted
  signal incrementNumberOfPacketsTransmitted_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal incrementNumberOfPacketsTransmitted_tag_out   : std_logic_vector(1 downto 0);
  signal incrementNumberOfPacketsTransmitted_start_req : std_logic;
  signal incrementNumberOfPacketsTransmitted_start_ack : std_logic;
  signal incrementNumberOfPacketsTransmitted_fin_req   : std_logic;
  signal incrementNumberOfPacketsTransmitted_fin_ack : std_logic;
  -- caller side aggregated signals for module incrementNumberOfPacketsTransmitted
  signal incrementNumberOfPacketsTransmitted_call_reqs: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsTransmitted_call_acks: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsTransmitted_return_reqs: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsTransmitted_return_acks: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsTransmitted_call_tag: std_logic_vector(0 downto 0);
  signal incrementNumberOfPacketsTransmitted_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module incrementRegister
  component incrementRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      reg_index : in  std_logic_vector(7 downto 0);
      incremented_value : out  std_logic_vector(31 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module incrementRegister
  signal incrementRegister_reg_index :  std_logic_vector(7 downto 0);
  signal incrementRegister_incremented_value :  std_logic_vector(31 downto 0);
  signal incrementRegister_in_args    : std_logic_vector(7 downto 0);
  signal incrementRegister_out_args   : std_logic_vector(31 downto 0);
  signal incrementRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal incrementRegister_tag_out   : std_logic_vector(2 downto 0);
  signal incrementRegister_start_req : std_logic;
  signal incrementRegister_start_ack : std_logic;
  signal incrementRegister_fin_req   : std_logic;
  signal incrementRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module incrementRegister
  signal incrementRegister_call_reqs: std_logic_vector(1 downto 0);
  signal incrementRegister_call_acks: std_logic_vector(1 downto 0);
  signal incrementRegister_return_reqs: std_logic_vector(1 downto 0);
  signal incrementRegister_return_acks: std_logic_vector(1 downto 0);
  signal incrementRegister_call_data: std_logic_vector(15 downto 0);
  signal incrementRegister_call_tag: std_logic_vector(1 downto 0);
  signal incrementRegister_return_data: std_logic_vector(63 downto 0);
  signal incrementRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      max_addr_offset : in  std_logic_vector(15 downto 0);
      rx_buffer_pointer : in  std_logic_vector(63 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(71 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(15 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(103 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(106 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_tag :  std_logic_vector(7 downto 0);
  signal loadBuffer_max_addr_offset :  std_logic_vector(15 downto 0);
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(63 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(87 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(87 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      S_CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(1 downto 0);
      accessRegister_call_acks : in   std_logic_vector(1 downto 0);
      accessRegister_call_data : out  std_logic_vector(89 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(1 downto 0);
      accessRegister_return_acks : in   std_logic_vector(1 downto 0);
      accessRegister_return_data : in   std_logic_vector(63 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_r_data : out  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueMisc_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueMisc_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueMisc_call_data : out  std_logic_vector(104 downto 0);
      accessQueueMisc_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueMisc_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueMisc_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueMisc_return_data : in   std_logic_vector(31 downto 0);
      accessQueueMisc_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(103 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(63 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_tag :  std_logic_vector(7 downto 0);
  signal popFromQueue_queue_type :  std_logic_vector(1 downto 0);
  signal popFromQueue_server_id :  std_logic_vector(7 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(63 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(17 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(64 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(35 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(129 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      rx_buffer_pointer : in  std_logic_vector(63 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(7 downto 0);
      S_NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(7 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_call_reqs : out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_call_acks : in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_return_reqs : out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_return_acks : in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsReceived_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_tag :  std_logic_vector(7 downto 0);
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(63 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(71 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(71 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      queue_type : in  std_logic_vector(1 downto 0);
      server_id : in  std_logic_vector(7 downto 0);
      q_w_data : in  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_req : out  std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_ack : in   std_logic_vector(0 downto 0);
      QUEUE_MONITOR_SIGNAL_pipe_write_data : out  std_logic_vector(31 downto 0);
      getQueuePointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_call_data : out  std_logic_vector(9 downto 0);
      getQueuePointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointer_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointer_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueLockPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLockPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLockPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueLockPointer_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_call_data : out  std_logic_vector(168 downto 0);
      accessMemoryWord_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryWord_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryWord_return_data : in   std_logic_vector(31 downto 0);
      accessMemoryWord_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(71 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      setTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_call_data : out  std_logic_vector(103 downto 0);
      setTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      setTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      setTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      setTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(135 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(71 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(71 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_call_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_call_data : out  std_logic_vector(9 downto 0);
      getQueueBufPointer_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueBufPointer_return_acks : in   std_logic_vector(0 downto 0);
      getQueueBufPointer_return_data : in   std_logic_vector(63 downto 0);
      getQueueBufPointer_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(71 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(71 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(167 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_tag :  std_logic_vector(7 downto 0);
  signal pushIntoQueue_queue_type :  std_logic_vector(1 downto 0);
  signal pushIntoQueue_server_id :  std_logic_vector(7 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(63 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(81 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(245 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseLock
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      lock_address_pointer : in  std_logic_vector(63 downto 0);
      accessMemoryByte_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByte_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByte_call_data : out  std_logic_vector(144 downto 0);
      accessMemoryByte_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMemoryByte_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryByte_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryByte_return_data : in   std_logic_vector(7 downto 0);
      accessMemoryByte_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseLock
  signal releaseLock_tag :  std_logic_vector(7 downto 0);
  signal releaseLock_lock_address_pointer :  std_logic_vector(63 downto 0);
  signal releaseLock_in_args    : std_logic_vector(71 downto 0);
  signal releaseLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseLock_tag_out   : std_logic_vector(2 downto 0);
  signal releaseLock_start_req : std_logic;
  signal releaseLock_start_ack : std_logic;
  signal releaseLock_fin_req   : std_logic;
  signal releaseLock_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseLock
  signal releaseLock_call_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_call_acks: std_logic_vector(1 downto 0);
  signal releaseLock_return_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_return_acks: std_logic_vector(1 downto 0);
  signal releaseLock_call_data: std_logic_vector(143 downto 0);
  signal releaseLock_call_tag: std_logic_vector(1 downto 0);
  signal releaseLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setGlobalSignals
  component setGlobalSignals is -- 
    generic (tag_length : integer); 
    port ( -- 
      NIC_INTR_ENABLE : in std_logic_vector(0 downto 0);
      NIC_INTR_INTERNAL : in std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_pipe_write_data : out  std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_INTR_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      S_CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      S_NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      accessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_call_acks : in   std_logic_vector(0 downto 0);
      accessRegister_call_data : out  std_logic_vector(44 downto 0);
      accessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      accessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      accessRegister_return_acks : in   std_logic_vector(0 downto 0);
      accessRegister_return_data : in   std_logic_vector(31 downto 0);
      accessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setGlobalSignals
  signal setGlobalSignals_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setGlobalSignals_tag_out   : std_logic_vector(1 downto 0);
  signal setGlobalSignals_start_req : std_logic;
  signal setGlobalSignals_start_ack : std_logic;
  signal setGlobalSignals_fin_req   : std_logic;
  signal setGlobalSignals_fin_ack : std_logic;
  -- caller side aggregated signals for module setGlobalSignals
  signal setGlobalSignals_call_reqs: std_logic_vector(0 downto 0);
  signal setGlobalSignals_call_acks: std_logic_vector(0 downto 0);
  signal setGlobalSignals_return_reqs: std_logic_vector(0 downto 0);
  signal setGlobalSignals_return_acks: std_logic_vector(0 downto 0);
  signal setGlobalSignals_call_tag: std_logic_vector(0 downto 0);
  signal setGlobalSignals_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      buf_base_address : in  std_logic_vector(63 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(63 downto 0);
      accessQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_call_data : out  std_logic_vector(168 downto 0);
      accessQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueElement_return_data : in   std_logic_vector(63 downto 0);
      accessQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_tag :  std_logic_vector(7 downto 0);
  signal setQueueElement_buf_base_address :  std_logic_vector(63 downto 0);
  signal setQueueElement_write_index :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(63 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(167 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(167 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessQueueReadIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueReadIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueReadIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueReadIndex_return_tag :  in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_call_data : out  std_logic_vector(104 downto 0);
      accessQueueWriteIndex_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueWriteIndex_return_data : in   std_logic_vector(31 downto 0);
      accessQueueWriteIndex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_tag :  std_logic_vector(7 downto 0);
  signal setQueuePointers_q_base_address :  std_logic_vector(63 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(135 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(271 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setTotalMessages
  component setTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      q_base_address : in  std_logic_vector(63 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_call_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_call_data : out  std_logic_vector(104 downto 0);
      accessQueueTotalMsgs_call_tag  :  out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_reqs : out  std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_acks : in   std_logic_vector(0 downto 0);
      accessQueueTotalMsgs_return_data : in   std_logic_vector(31 downto 0);
      accessQueueTotalMsgs_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setTotalMessages
  signal setTotalMessages_tag :  std_logic_vector(7 downto 0);
  signal setTotalMessages_q_base_address :  std_logic_vector(63 downto 0);
  signal setTotalMessages_updated_total_msgs :  std_logic_vector(31 downto 0);
  signal setTotalMessages_in_args    : std_logic_vector(103 downto 0);
  signal setTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal setTotalMessages_start_req : std_logic;
  signal setTotalMessages_start_ack : std_logic;
  signal setTotalMessages_fin_req   : std_logic;
  signal setTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module setTotalMessages
  signal setTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal setTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal setTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal setTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal setTotalMessages_call_data: std_logic_vector(207 downto 0);
  signal setTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal setTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(7 downto 0);
      S_CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      S_NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(15 downto 0);
      TX_ACTIVITY_LOGGER_pipe_write_req : out  std_logic_vector(0 downto 0);
      TX_ACTIVITY_LOGGER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      TX_ACTIVITY_LOGGER_pipe_write_data : out  std_logic_vector(7 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(81 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(15 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(64 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsTransmitted_call_reqs : out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsTransmitted_call_acks : in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsTransmitted_call_tag  :  out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsTransmitted_return_reqs : out  std_logic_vector(0 downto 0);
      incrementNumberOfPacketsTransmitted_return_acks : in   std_logic_vector(0 downto 0);
      incrementNumberOfPacketsTransmitted_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(71 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      packet_pointer : in  std_logic_vector(63 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(1 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(401 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(1 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(127 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_tag :  std_logic_vector(7 downto 0);
  signal transmitPacket_packet_pointer :  std_logic_vector(63 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(71 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(71 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      base_buffer_pointer : in  std_logic_vector(63 downto 0);
      max_addr_offset : in  std_logic_vector(15 downto 0);
      packet_size : in  std_logic_vector(10 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_tag :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(63 downto 0);
  signal writeControlInformationToMem_max_addr_offset :  std_logic_vector(15 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(10 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(106 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(106 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      buf_pointer : in  std_logic_vector(63 downto 0);
      addr_offset : out  std_logic_vector(15 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_tag :  std_logic_vector(7 downto 0);
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(63 downto 0);
  signal writeEthernetHeaderToMem_addr_offset :  std_logic_vector(15 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(71 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(15 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(71 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(15 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      tag : in  std_logic_vector(7 downto 0);
      max_addr_offset : in  std_logic_vector(15 downto 0);
      base_buf_pointer : in  std_logic_vector(63 downto 0);
      addr_offset : in  std_logic_vector(15 downto 0);
      packet_size_11 : out  std_logic_vector(10 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemoryDword_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_call_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_call_data : out  std_logic_vector(200 downto 0);
      accessMemoryDword_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemoryDword_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemoryDword_return_acks : in   std_logic_vector(0 downto 0);
      accessMemoryDword_return_data : in   std_logic_vector(63 downto 0);
      accessMemoryDword_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_tag :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_max_addr_offset :  std_logic_vector(15 downto 0);
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(63 downto 0);
  signal writePayloadToMem_addr_offset :  std_logic_vector(15 downto 0);
  signal writePayloadToMem_packet_size_11 :  std_logic_vector(10 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(103 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(19 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(103 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(19 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(15 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(7 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(15 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(7 downto 0);
  -- aggregate signals for write to pipe MAC_ENABLE
  signal MAC_ENABLE_pipe_write_data: std_logic_vector(1 downto 0);
  signal MAC_ENABLE_pipe_write_req: std_logic_vector(1 downto 0);
  signal MAC_ENABLE_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_DEBUG_SIGNAL
  signal NIC_DEBUG_SIGNAL_pipe_write_data: std_logic_vector(255 downto 0);
  signal NIC_DEBUG_SIGNAL_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_DEBUG_SIGNAL_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_INTR
  signal NIC_INTR_pipe_write_data: std_logic_vector(1 downto 0);
  signal NIC_INTR_pipe_write_req: std_logic_vector(1 downto 0);
  signal NIC_INTR_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe NIC_INTR_ENABLE
  signal NIC_INTR_ENABLE_pipe_write_data: std_logic_vector(1 downto 0);
  signal NIC_INTR_ENABLE_pipe_write_req: std_logic_vector(1 downto 0);
  signal NIC_INTR_ENABLE_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe NIC_INTR_ENABLE
  signal NIC_INTR_ENABLE: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_INTR_INTERNAL
  signal NIC_INTR_INTERNAL_pipe_write_data: std_logic_vector(0 downto 0);
  signal NIC_INTR_INTERNAL_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_INTR_INTERNAL_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NIC_INTR_INTERNAL
  signal NIC_INTR_INTERNAL: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe QUEUE_MONITOR_SIGNAL
  signal QUEUE_MONITOR_SIGNAL_pipe_write_data: std_logic_vector(63 downto 0);
  signal QUEUE_MONITOR_SIGNAL_pipe_write_req: std_logic_vector(1 downto 0);
  signal QUEUE_MONITOR_SIGNAL_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe QUEUE_MONITOR_SIGNAL
  signal QUEUE_MONITOR_SIGNAL: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe RX_ACTIVITY_LOGGER
  signal RX_ACTIVITY_LOGGER_pipe_write_data: std_logic_vector(7 downto 0);
  signal RX_ACTIVITY_LOGGER_pipe_write_req: std_logic_vector(0 downto 0);
  signal RX_ACTIVITY_LOGGER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe S_CONTROL_REGISTER
  signal S_CONTROL_REGISTER_pipe_write_data: std_logic_vector(63 downto 0);
  signal S_CONTROL_REGISTER_pipe_write_req: std_logic_vector(1 downto 0);
  signal S_CONTROL_REGISTER_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe S_CONTROL_REGISTER
  signal S_CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe S_NUMBER_OF_SERVERS
  signal S_NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(63 downto 0);
  signal S_NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(1 downto 0);
  signal S_NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe S_NUMBER_OF_SERVERS
  signal S_NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe TX_ACTIVITY_LOGGER
  signal TX_ACTIVITY_LOGGER_pipe_write_data: std_logic_vector(7 downto 0);
  signal TX_ACTIVITY_LOGGER_pipe_write_req: std_logic_vector(0 downto 0);
  signal TX_ACTIVITY_LOGGER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe memory_access_lock
  signal memory_access_lock_pipe_write_data: std_logic_vector(1 downto 0);
  signal memory_access_lock_pipe_write_req: std_logic_vector(1 downto 0);
  signal memory_access_lock_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe memory_access_lock
  signal memory_access_lock_pipe_read_data: std_logic_vector(0 downto 0);
  signal memory_access_lock_pipe_read_req: std_logic_vector(0 downto 0);
  signal memory_access_lock_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(145 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      S_CONTROL_REGISTER => S_CONTROL_REGISTER,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(7 downto 0),
      RX_ACTIVITY_LOGGER_pipe_write_req => RX_ACTIVITY_LOGGER_pipe_write_req(0 downto 0),
      RX_ACTIVITY_LOGGER_pipe_write_ack => RX_ACTIVITY_LOGGER_pipe_write_ack(0 downto 0),
      RX_ACTIVITY_LOGGER_pipe_write_data => RX_ACTIVITY_LOGGER_pipe_write_data(7 downto 0),
      accessRegister_call_reqs => accessRegister_call_reqs(5 downto 5),
      accessRegister_call_acks => accessRegister_call_acks(5 downto 5),
      accessRegister_call_data => accessRegister_call_data(269 downto 225),
      accessRegister_call_tag => accessRegister_call_tag(11 downto 10),
      accessRegister_return_reqs => accessRegister_return_reqs(5 downto 5),
      accessRegister_return_acks => accessRegister_return_acks(5 downto 5),
      accessRegister_return_data => accessRegister_return_data(191 downto 160),
      accessRegister_return_tag => accessRegister_return_tag(11 downto 10),
      accessMemoryDword_call_reqs => accessMemoryDword_call_reqs(2 downto 2),
      accessMemoryDword_call_acks => accessMemoryDword_call_acks(2 downto 2),
      accessMemoryDword_call_data => accessMemoryDword_call_data(602 downto 402),
      accessMemoryDword_call_tag => accessMemoryDword_call_tag(5 downto 4),
      accessMemoryDword_return_reqs => accessMemoryDword_return_reqs(2 downto 2),
      accessMemoryDword_return_acks => accessMemoryDword_return_acks(2 downto 2),
      accessMemoryDword_return_data => accessMemoryDword_return_data(191 downto 128),
      accessMemoryDword_return_tag => accessMemoryDword_return_tag(5 downto 4),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(35 downto 18),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(129 downto 65),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(87 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(163 downto 82),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(71 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module accessMemoryBase
  accessMemoryBase_tag <= accessMemoryBase_in_args(117 downto 110);
  accessMemoryBase_request <= accessMemoryBase_in_args(109 downto 0);
  accessMemoryBase_out_args <= accessMemoryBase_response ;
  -- call arbiter for module accessMemoryBase
  accessMemoryBase_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 118,
      return_data_width => 65,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMemoryBase_call_reqs,
      call_acks => accessMemoryBase_call_acks,
      return_reqs => accessMemoryBase_return_reqs,
      return_acks => accessMemoryBase_return_acks,
      call_data  => accessMemoryBase_call_data,
      call_tag  => accessMemoryBase_call_tag,
      return_tag  => accessMemoryBase_return_tag,
      call_mtag => accessMemoryBase_tag_in,
      return_mtag => accessMemoryBase_tag_out,
      return_data =>accessMemoryBase_return_data,
      call_mreq => accessMemoryBase_start_req,
      call_mack => accessMemoryBase_start_ack,
      return_mreq => accessMemoryBase_fin_req,
      return_mack => accessMemoryBase_fin_ack,
      call_mdata => accessMemoryBase_in_args,
      return_mdata => accessMemoryBase_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryBase_instance:accessMemoryBase-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => accessMemoryBase_tag,
      request => accessMemoryBase_request,
      response => accessMemoryBase_response,
      start_req => accessMemoryBase_start_req,
      start_ack => accessMemoryBase_start_ack,
      fin_req => accessMemoryBase_fin_req,
      fin_ack => accessMemoryBase_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_DEBUG_SIGNAL_pipe_write_req => NIC_DEBUG_SIGNAL_pipe_write_req(0 downto 0),
      NIC_DEBUG_SIGNAL_pipe_write_ack => NIC_DEBUG_SIGNAL_pipe_write_ack(0 downto 0),
      NIC_DEBUG_SIGNAL_pipe_write_data => NIC_DEBUG_SIGNAL_pipe_write_data(255 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemoryBase_tag_in,
      tag_out => accessMemoryBase_tag_out-- 
    ); -- 
  -- module accessMemoryByte
  accessMemoryByte_tag <= accessMemoryByte_in_args(144 downto 137);
  accessMemoryByte_rwbar <= accessMemoryByte_in_args(136 downto 136);
  accessMemoryByte_byte_addr_base <= accessMemoryByte_in_args(135 downto 72);
  accessMemoryByte_offset <= accessMemoryByte_in_args(71 downto 8);
  accessMemoryByte_wbyte <= accessMemoryByte_in_args(7 downto 0);
  accessMemoryByte_out_args <= accessMemoryByte_rbyte ;
  -- call arbiter for module accessMemoryByte
  accessMemoryByte_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 145,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMemoryByte_call_reqs,
      call_acks => accessMemoryByte_call_acks,
      return_reqs => accessMemoryByte_return_reqs,
      return_acks => accessMemoryByte_return_acks,
      call_data  => accessMemoryByte_call_data,
      call_tag  => accessMemoryByte_call_tag,
      return_tag  => accessMemoryByte_return_tag,
      call_mtag => accessMemoryByte_tag_in,
      return_mtag => accessMemoryByte_tag_out,
      return_data =>accessMemoryByte_return_data,
      call_mreq => accessMemoryByte_start_req,
      call_mack => accessMemoryByte_start_ack,
      return_mreq => accessMemoryByte_fin_req,
      return_mack => accessMemoryByte_fin_ack,
      call_mdata => accessMemoryByte_in_args,
      return_mdata => accessMemoryByte_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryByte_instance:accessMemoryByte-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => accessMemoryByte_tag,
      rwbar => accessMemoryByte_rwbar,
      byte_addr_base => accessMemoryByte_byte_addr_base,
      offset => accessMemoryByte_offset,
      wbyte => accessMemoryByte_wbyte,
      rbyte => accessMemoryByte_rbyte,
      start_req => accessMemoryByte_start_req,
      start_ack => accessMemoryByte_start_ack,
      fin_req => accessMemoryByte_fin_req,
      fin_ack => accessMemoryByte_fin_ack,
      clk => clk,
      reset => reset,
      doMemAccess_call_reqs => doMemAccess_call_reqs(1 downto 1),
      doMemAccess_call_acks => doMemAccess_call_acks(1 downto 1),
      doMemAccess_call_data => doMemAccess_call_data(405 downto 203),
      doMemAccess_call_tag => doMemAccess_call_tag(1 downto 1),
      doMemAccess_return_reqs => doMemAccess_return_reqs(1 downto 1),
      doMemAccess_return_acks => doMemAccess_return_acks(1 downto 1),
      doMemAccess_return_data => doMemAccess_return_data(127 downto 64),
      doMemAccess_return_tag => doMemAccess_return_tag(1 downto 1),
      tag_in => accessMemoryByte_tag_in,
      tag_out => accessMemoryByte_tag_out-- 
    ); -- 
  -- module accessMemoryByteBase
  accessMemoryByteBase_tag <= accessMemoryByteBase_in_args(145 downto 138);
  accessMemoryByteBase_lock <= accessMemoryByteBase_in_args(137 downto 137);
  accessMemoryByteBase_rwbar <= accessMemoryByteBase_in_args(136 downto 136);
  accessMemoryByteBase_byte_addr_base <= accessMemoryByteBase_in_args(135 downto 72);
  accessMemoryByteBase_offset <= accessMemoryByteBase_in_args(71 downto 8);
  accessMemoryByteBase_wbyte <= accessMemoryByteBase_in_args(7 downto 0);
  accessMemoryByteBase_out_args <= accessMemoryByteBase_rbyte ;
  -- call arbiter for module accessMemoryByteBase
  accessMemoryByteBase_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 146,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMemoryByteBase_call_reqs,
      call_acks => accessMemoryByteBase_call_acks,
      return_reqs => accessMemoryByteBase_return_reqs,
      return_acks => accessMemoryByteBase_return_acks,
      call_data  => accessMemoryByteBase_call_data,
      call_tag  => accessMemoryByteBase_call_tag,
      return_tag  => accessMemoryByteBase_return_tag,
      call_mtag => accessMemoryByteBase_tag_in,
      return_mtag => accessMemoryByteBase_tag_out,
      return_data =>accessMemoryByteBase_return_data,
      call_mreq => accessMemoryByteBase_start_req,
      call_mack => accessMemoryByteBase_start_ack,
      return_mreq => accessMemoryByteBase_fin_req,
      return_mack => accessMemoryByteBase_fin_ack,
      call_mdata => accessMemoryByteBase_in_args,
      return_mdata => accessMemoryByteBase_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryByteBase_instance:accessMemoryByteBase-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => accessMemoryByteBase_tag,
      lock => accessMemoryByteBase_lock,
      rwbar => accessMemoryByteBase_rwbar,
      byte_addr_base => accessMemoryByteBase_byte_addr_base,
      offset => accessMemoryByteBase_offset,
      wbyte => accessMemoryByteBase_wbyte,
      rbyte => accessMemoryByteBase_rbyte,
      start_req => accessMemoryByteBase_start_req,
      start_ack => accessMemoryByteBase_start_ack,
      fin_req => accessMemoryByteBase_fin_req,
      fin_ack => accessMemoryByteBase_fin_ack,
      clk => clk,
      reset => reset,
      calculateAddress36_call_reqs => calculateAddress36_call_reqs(1 downto 1),
      calculateAddress36_call_acks => calculateAddress36_call_acks(1 downto 1),
      calculateAddress36_call_data => calculateAddress36_call_data(255 downto 128),
      calculateAddress36_call_tag => calculateAddress36_call_tag(1 downto 1),
      calculateAddress36_return_reqs => calculateAddress36_return_reqs(1 downto 1),
      calculateAddress36_return_acks => calculateAddress36_return_acks(1 downto 1),
      calculateAddress36_return_data => calculateAddress36_return_data(71 downto 36),
      calculateAddress36_return_tag => calculateAddress36_return_tag(1 downto 1),
      accessMemoryBase_call_reqs => accessMemoryBase_call_reqs(1 downto 1),
      accessMemoryBase_call_acks => accessMemoryBase_call_acks(1 downto 1),
      accessMemoryBase_call_data => accessMemoryBase_call_data(235 downto 118),
      accessMemoryBase_call_tag => accessMemoryBase_call_tag(1 downto 1),
      accessMemoryBase_return_reqs => accessMemoryBase_return_reqs(1 downto 1),
      accessMemoryBase_return_acks => accessMemoryBase_return_acks(1 downto 1),
      accessMemoryBase_return_data => accessMemoryBase_return_data(129 downto 65),
      accessMemoryBase_return_tag => accessMemoryBase_return_tag(1 downto 1),
      tag_in => accessMemoryByteBase_tag_in,
      tag_out => accessMemoryByteBase_tag_out-- 
    ); -- 
  -- module accessMemoryDword
  accessMemoryDword_tag <= accessMemoryDword_in_args(200 downto 193);
  accessMemoryDword_rwbar <= accessMemoryDword_in_args(192 downto 192);
  accessMemoryDword_base_addr <= accessMemoryDword_in_args(191 downto 128);
  accessMemoryDword_offset <= accessMemoryDword_in_args(127 downto 64);
  accessMemoryDword_wdata <= accessMemoryDword_in_args(63 downto 0);
  accessMemoryDword_out_args <= accessMemoryDword_rdata ;
  -- call arbiter for module accessMemoryDword
  accessMemoryDword_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 7,
      call_data_width => 201,
      return_data_width => 64,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMemoryDword_call_reqs,
      call_acks => accessMemoryDword_call_acks,
      return_reqs => accessMemoryDword_return_reqs,
      return_acks => accessMemoryDword_return_acks,
      call_data  => accessMemoryDword_call_data,
      call_tag  => accessMemoryDword_call_tag,
      return_tag  => accessMemoryDword_return_tag,
      call_mtag => accessMemoryDword_tag_in,
      return_mtag => accessMemoryDword_tag_out,
      return_data =>accessMemoryDword_return_data,
      call_mreq => accessMemoryDword_start_req,
      call_mack => accessMemoryDword_start_ack,
      return_mreq => accessMemoryDword_fin_req,
      return_mack => accessMemoryDword_fin_ack,
      call_mdata => accessMemoryDword_in_args,
      return_mdata => accessMemoryDword_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryDword_instance:accessMemoryDword-- 
    generic map(tag_length => 5)
    port map(-- 
      tag => accessMemoryDword_tag,
      rwbar => accessMemoryDword_rwbar,
      base_addr => accessMemoryDword_base_addr,
      offset => accessMemoryDword_offset,
      wdata => accessMemoryDword_wdata,
      rdata => accessMemoryDword_rdata,
      start_req => accessMemoryDword_start_req,
      start_ack => accessMemoryDword_start_ack,
      fin_req => accessMemoryDword_fin_req,
      fin_ack => accessMemoryDword_fin_ack,
      clk => clk,
      reset => reset,
      doMemAccess_call_reqs => doMemAccess_call_reqs(0 downto 0),
      doMemAccess_call_acks => doMemAccess_call_acks(0 downto 0),
      doMemAccess_call_data => doMemAccess_call_data(202 downto 0),
      doMemAccess_call_tag => doMemAccess_call_tag(0 downto 0),
      doMemAccess_return_reqs => doMemAccess_return_reqs(0 downto 0),
      doMemAccess_return_acks => doMemAccess_return_acks(0 downto 0),
      doMemAccess_return_data => doMemAccess_return_data(63 downto 0),
      doMemAccess_return_tag => doMemAccess_return_tag(0 downto 0),
      tag_in => accessMemoryDword_tag_in,
      tag_out => accessMemoryDword_tag_out-- 
    ); -- 
  -- module accessMemoryDwordBase
  accessMemoryDwordBase_tag <= accessMemoryDwordBase_in_args(201 downto 194);
  accessMemoryDwordBase_lock <= accessMemoryDwordBase_in_args(193 downto 193);
  accessMemoryDwordBase_rwbar <= accessMemoryDwordBase_in_args(192 downto 192);
  accessMemoryDwordBase_base_addr <= accessMemoryDwordBase_in_args(191 downto 128);
  accessMemoryDwordBase_offset <= accessMemoryDwordBase_in_args(127 downto 64);
  accessMemoryDwordBase_wdata <= accessMemoryDwordBase_in_args(63 downto 0);
  accessMemoryDwordBase_out_args <= accessMemoryDwordBase_rdata ;
  -- call arbiter for module accessMemoryDwordBase
  accessMemoryDwordBase_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 202,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMemoryDwordBase_call_reqs,
      call_acks => accessMemoryDwordBase_call_acks,
      return_reqs => accessMemoryDwordBase_return_reqs,
      return_acks => accessMemoryDwordBase_return_acks,
      call_data  => accessMemoryDwordBase_call_data,
      call_tag  => accessMemoryDwordBase_call_tag,
      return_tag  => accessMemoryDwordBase_return_tag,
      call_mtag => accessMemoryDwordBase_tag_in,
      return_mtag => accessMemoryDwordBase_tag_out,
      return_data =>accessMemoryDwordBase_return_data,
      call_mreq => accessMemoryDwordBase_start_req,
      call_mack => accessMemoryDwordBase_start_ack,
      return_mreq => accessMemoryDwordBase_fin_req,
      return_mack => accessMemoryDwordBase_fin_ack,
      call_mdata => accessMemoryDwordBase_in_args,
      return_mdata => accessMemoryDwordBase_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryDwordBase_instance:accessMemoryDwordBase-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => accessMemoryDwordBase_tag,
      lock => accessMemoryDwordBase_lock,
      rwbar => accessMemoryDwordBase_rwbar,
      base_addr => accessMemoryDwordBase_base_addr,
      offset => accessMemoryDwordBase_offset,
      wdata => accessMemoryDwordBase_wdata,
      rdata => accessMemoryDwordBase_rdata,
      start_req => accessMemoryDwordBase_start_req,
      start_ack => accessMemoryDwordBase_start_ack,
      fin_req => accessMemoryDwordBase_fin_req,
      fin_ack => accessMemoryDwordBase_fin_ack,
      clk => clk,
      reset => reset,
      calculateAddress36_call_reqs => calculateAddress36_call_reqs(0 downto 0),
      calculateAddress36_call_acks => calculateAddress36_call_acks(0 downto 0),
      calculateAddress36_call_data => calculateAddress36_call_data(127 downto 0),
      calculateAddress36_call_tag => calculateAddress36_call_tag(0 downto 0),
      calculateAddress36_return_reqs => calculateAddress36_return_reqs(0 downto 0),
      calculateAddress36_return_acks => calculateAddress36_return_acks(0 downto 0),
      calculateAddress36_return_data => calculateAddress36_return_data(35 downto 0),
      calculateAddress36_return_tag => calculateAddress36_return_tag(0 downto 0),
      accessMemoryBase_call_reqs => accessMemoryBase_call_reqs(0 downto 0),
      accessMemoryBase_call_acks => accessMemoryBase_call_acks(0 downto 0),
      accessMemoryBase_call_data => accessMemoryBase_call_data(117 downto 0),
      accessMemoryBase_call_tag => accessMemoryBase_call_tag(0 downto 0),
      accessMemoryBase_return_reqs => accessMemoryBase_return_reqs(0 downto 0),
      accessMemoryBase_return_acks => accessMemoryBase_return_acks(0 downto 0),
      accessMemoryBase_return_data => accessMemoryBase_return_data(64 downto 0),
      accessMemoryBase_return_tag => accessMemoryBase_return_tag(0 downto 0),
      tag_in => accessMemoryDwordBase_tag_in,
      tag_out => accessMemoryDwordBase_tag_out-- 
    ); -- 
  -- module accessMemoryLdStub
  accessMemoryLdStub_tag <= accessMemoryLdStub_in_args(135 downto 128);
  accessMemoryLdStub_byte_addr_base <= accessMemoryLdStub_in_args(127 downto 64);
  accessMemoryLdStub_offset <= accessMemoryLdStub_in_args(63 downto 0);
  accessMemoryLdStub_out_args <= accessMemoryLdStub_rbyte ;
  -- call arbiter for module accessMemoryLdStub
  accessMemoryLdStub_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 136,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMemoryLdStub_call_reqs,
      call_acks => accessMemoryLdStub_call_acks,
      return_reqs => accessMemoryLdStub_return_reqs,
      return_acks => accessMemoryLdStub_return_acks,
      call_data  => accessMemoryLdStub_call_data,
      call_tag  => accessMemoryLdStub_call_tag,
      return_tag  => accessMemoryLdStub_return_tag,
      call_mtag => accessMemoryLdStub_tag_in,
      return_mtag => accessMemoryLdStub_tag_out,
      return_data =>accessMemoryLdStub_return_data,
      call_mreq => accessMemoryLdStub_start_req,
      call_mack => accessMemoryLdStub_start_ack,
      return_mreq => accessMemoryLdStub_fin_req,
      return_mack => accessMemoryLdStub_fin_ack,
      call_mdata => accessMemoryLdStub_in_args,
      return_mdata => accessMemoryLdStub_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryLdStub_instance:accessMemoryLdStub-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => accessMemoryLdStub_tag,
      byte_addr_base => accessMemoryLdStub_byte_addr_base,
      offset => accessMemoryLdStub_offset,
      rbyte => accessMemoryLdStub_rbyte,
      start_req => accessMemoryLdStub_start_req,
      start_ack => accessMemoryLdStub_start_ack,
      fin_req => accessMemoryLdStub_fin_req,
      fin_ack => accessMemoryLdStub_fin_ack,
      clk => clk,
      reset => reset,
      doMemAccess_call_reqs => doMemAccess_call_reqs(3 downto 3),
      doMemAccess_call_acks => doMemAccess_call_acks(3 downto 3),
      doMemAccess_call_data => doMemAccess_call_data(811 downto 609),
      doMemAccess_call_tag => doMemAccess_call_tag(3 downto 3),
      doMemAccess_return_reqs => doMemAccess_return_reqs(3 downto 3),
      doMemAccess_return_acks => doMemAccess_return_acks(3 downto 3),
      doMemAccess_return_data => doMemAccess_return_data(255 downto 192),
      doMemAccess_return_tag => doMemAccess_return_tag(3 downto 3),
      tag_in => accessMemoryLdStub_tag_in,
      tag_out => accessMemoryLdStub_tag_out-- 
    ); -- 
  -- module accessMemoryWord
  accessMemoryWord_tag <= accessMemoryWord_in_args(168 downto 161);
  accessMemoryWord_rwbar <= accessMemoryWord_in_args(160 downto 160);
  accessMemoryWord_word_addr_base <= accessMemoryWord_in_args(159 downto 96);
  accessMemoryWord_offset <= accessMemoryWord_in_args(95 downto 32);
  accessMemoryWord_wword <= accessMemoryWord_in_args(31 downto 0);
  accessMemoryWord_out_args <= accessMemoryWord_rword ;
  -- call arbiter for module accessMemoryWord
  accessMemoryWord_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 6,
      call_data_width => 169,
      return_data_width => 32,
      callee_tag_length => 3,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMemoryWord_call_reqs,
      call_acks => accessMemoryWord_call_acks,
      return_reqs => accessMemoryWord_return_reqs,
      return_acks => accessMemoryWord_return_acks,
      call_data  => accessMemoryWord_call_data,
      call_tag  => accessMemoryWord_call_tag,
      return_tag  => accessMemoryWord_return_tag,
      call_mtag => accessMemoryWord_tag_in,
      return_mtag => accessMemoryWord_tag_out,
      return_data =>accessMemoryWord_return_data,
      call_mreq => accessMemoryWord_start_req,
      call_mack => accessMemoryWord_start_ack,
      return_mreq => accessMemoryWord_fin_req,
      return_mack => accessMemoryWord_fin_ack,
      call_mdata => accessMemoryWord_in_args,
      return_mdata => accessMemoryWord_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryWord_instance:accessMemoryWord-- 
    generic map(tag_length => 4)
    port map(-- 
      tag => accessMemoryWord_tag,
      rwbar => accessMemoryWord_rwbar,
      word_addr_base => accessMemoryWord_word_addr_base,
      offset => accessMemoryWord_offset,
      wword => accessMemoryWord_wword,
      rword => accessMemoryWord_rword,
      start_req => accessMemoryWord_start_req,
      start_ack => accessMemoryWord_start_ack,
      fin_req => accessMemoryWord_fin_req,
      fin_ack => accessMemoryWord_fin_ack,
      clk => clk,
      reset => reset,
      doMemAccess_call_reqs => doMemAccess_call_reqs(2 downto 2),
      doMemAccess_call_acks => doMemAccess_call_acks(2 downto 2),
      doMemAccess_call_data => doMemAccess_call_data(608 downto 406),
      doMemAccess_call_tag => doMemAccess_call_tag(2 downto 2),
      doMemAccess_return_reqs => doMemAccess_return_reqs(2 downto 2),
      doMemAccess_return_acks => doMemAccess_return_acks(2 downto 2),
      doMemAccess_return_data => doMemAccess_return_data(191 downto 128),
      doMemAccess_return_tag => doMemAccess_return_tag(2 downto 2),
      tag_in => accessMemoryWord_tag_in,
      tag_out => accessMemoryWord_tag_out-- 
    ); -- 
  -- module accessMemoryWordBase
  accessMemoryWordBase_tag <= accessMemoryWordBase_in_args(169 downto 162);
  accessMemoryWordBase_lock <= accessMemoryWordBase_in_args(161 downto 161);
  accessMemoryWordBase_rwbar <= accessMemoryWordBase_in_args(160 downto 160);
  accessMemoryWordBase_word_addr_base <= accessMemoryWordBase_in_args(159 downto 96);
  accessMemoryWordBase_offset <= accessMemoryWordBase_in_args(95 downto 32);
  accessMemoryWordBase_wword <= accessMemoryWordBase_in_args(31 downto 0);
  accessMemoryWordBase_out_args <= accessMemoryWordBase_rword ;
  -- call arbiter for module accessMemoryWordBase
  accessMemoryWordBase_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 170,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMemoryWordBase_call_reqs,
      call_acks => accessMemoryWordBase_call_acks,
      return_reqs => accessMemoryWordBase_return_reqs,
      return_acks => accessMemoryWordBase_return_acks,
      call_data  => accessMemoryWordBase_call_data,
      call_tag  => accessMemoryWordBase_call_tag,
      return_tag  => accessMemoryWordBase_return_tag,
      call_mtag => accessMemoryWordBase_tag_in,
      return_mtag => accessMemoryWordBase_tag_out,
      return_data =>accessMemoryWordBase_return_data,
      call_mreq => accessMemoryWordBase_start_req,
      call_mack => accessMemoryWordBase_start_ack,
      return_mreq => accessMemoryWordBase_fin_req,
      return_mack => accessMemoryWordBase_fin_ack,
      call_mdata => accessMemoryWordBase_in_args,
      return_mdata => accessMemoryWordBase_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemoryWordBase_instance:accessMemoryWordBase-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => accessMemoryWordBase_tag,
      lock => accessMemoryWordBase_lock,
      rwbar => accessMemoryWordBase_rwbar,
      word_addr_base => accessMemoryWordBase_word_addr_base,
      offset => accessMemoryWordBase_offset,
      wword => accessMemoryWordBase_wword,
      rword => accessMemoryWordBase_rword,
      start_req => accessMemoryWordBase_start_req,
      start_ack => accessMemoryWordBase_start_ack,
      fin_req => accessMemoryWordBase_fin_req,
      fin_ack => accessMemoryWordBase_fin_ack,
      clk => clk,
      reset => reset,
      calculateAddress36_call_reqs => calculateAddress36_call_reqs(2 downto 2),
      calculateAddress36_call_acks => calculateAddress36_call_acks(2 downto 2),
      calculateAddress36_call_data => calculateAddress36_call_data(383 downto 256),
      calculateAddress36_call_tag => calculateAddress36_call_tag(2 downto 2),
      calculateAddress36_return_reqs => calculateAddress36_return_reqs(2 downto 2),
      calculateAddress36_return_acks => calculateAddress36_return_acks(2 downto 2),
      calculateAddress36_return_data => calculateAddress36_return_data(107 downto 72),
      calculateAddress36_return_tag => calculateAddress36_return_tag(2 downto 2),
      accessMemoryBase_call_reqs => accessMemoryBase_call_reqs(2 downto 2),
      accessMemoryBase_call_acks => accessMemoryBase_call_acks(2 downto 2),
      accessMemoryBase_call_data => accessMemoryBase_call_data(353 downto 236),
      accessMemoryBase_call_tag => accessMemoryBase_call_tag(2 downto 2),
      accessMemoryBase_return_reqs => accessMemoryBase_return_reqs(2 downto 2),
      accessMemoryBase_return_acks => accessMemoryBase_return_acks(2 downto 2),
      accessMemoryBase_return_data => accessMemoryBase_return_data(194 downto 130),
      accessMemoryBase_return_tag => accessMemoryBase_return_tag(2 downto 2),
      tag_in => accessMemoryWordBase_tag_in,
      tag_out => accessMemoryWordBase_tag_out-- 
    ); -- 
  -- module accessQueueElement
  accessQueueElement_tag <= accessQueueElement_in_args(168 downto 161);
  accessQueueElement_rwbar <= accessQueueElement_in_args(160 downto 160);
  accessQueueElement_base_addr <= accessQueueElement_in_args(159 downto 96);
  accessQueueElement_index <= accessQueueElement_in_args(95 downto 64);
  accessQueueElement_wdata <= accessQueueElement_in_args(63 downto 0);
  accessQueueElement_out_args <= accessQueueElement_rdata ;
  -- call arbiter for module accessQueueElement
  accessQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 169,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessQueueElement_call_reqs,
      call_acks => accessQueueElement_call_acks,
      return_reqs => accessQueueElement_return_reqs,
      return_acks => accessQueueElement_return_acks,
      call_data  => accessQueueElement_call_data,
      call_tag  => accessQueueElement_call_tag,
      return_tag  => accessQueueElement_return_tag,
      call_mtag => accessQueueElement_tag_in,
      return_mtag => accessQueueElement_tag_out,
      return_data =>accessQueueElement_return_data,
      call_mreq => accessQueueElement_start_req,
      call_mack => accessQueueElement_start_ack,
      return_mreq => accessQueueElement_fin_req,
      return_mack => accessQueueElement_fin_ack,
      call_mdata => accessQueueElement_in_args,
      return_mdata => accessQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessQueueElement_instance:accessQueueElement-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => accessQueueElement_tag,
      rwbar => accessQueueElement_rwbar,
      base_addr => accessQueueElement_base_addr,
      index => accessQueueElement_index,
      wdata => accessQueueElement_wdata,
      rdata => accessQueueElement_rdata,
      start_req => accessQueueElement_start_req,
      start_ack => accessQueueElement_start_ack,
      fin_req => accessQueueElement_fin_req,
      fin_ack => accessQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryDword_call_reqs => accessMemoryDword_call_reqs(5 downto 5),
      accessMemoryDword_call_acks => accessMemoryDword_call_acks(5 downto 5),
      accessMemoryDword_call_data => accessMemoryDword_call_data(1205 downto 1005),
      accessMemoryDword_call_tag => accessMemoryDword_call_tag(11 downto 10),
      accessMemoryDword_return_reqs => accessMemoryDword_return_reqs(5 downto 5),
      accessMemoryDword_return_acks => accessMemoryDword_return_acks(5 downto 5),
      accessMemoryDword_return_data => accessMemoryDword_return_data(383 downto 320),
      accessMemoryDword_return_tag => accessMemoryDword_return_tag(11 downto 10),
      tag_in => accessQueueElement_tag_in,
      tag_out => accessQueueElement_tag_out-- 
    ); -- 
  -- module accessQueueLength
  accessQueueLength_tag <= accessQueueLength_in_args(104 downto 97);
  accessQueueLength_rwbar <= accessQueueLength_in_args(96 downto 96);
  accessQueueLength_qptr <= accessQueueLength_in_args(95 downto 32);
  accessQueueLength_wdata <= accessQueueLength_in_args(31 downto 0);
  accessQueueLength_out_args <= accessQueueLength_rdata ;
  -- call arbiter for module accessQueueLength
  accessQueueLength_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 105,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessQueueLength_call_reqs,
      call_acks => accessQueueLength_call_acks,
      return_reqs => accessQueueLength_return_reqs,
      return_acks => accessQueueLength_return_acks,
      call_data  => accessQueueLength_call_data,
      call_tag  => accessQueueLength_call_tag,
      return_tag  => accessQueueLength_return_tag,
      call_mtag => accessQueueLength_tag_in,
      return_mtag => accessQueueLength_tag_out,
      return_data =>accessQueueLength_return_data,
      call_mreq => accessQueueLength_start_req,
      call_mack => accessQueueLength_start_ack,
      return_mreq => accessQueueLength_fin_req,
      return_mack => accessQueueLength_fin_ack,
      call_mdata => accessQueueLength_in_args,
      return_mdata => accessQueueLength_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessQueueLength_instance:accessQueueLength-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => accessQueueLength_tag,
      rwbar => accessQueueLength_rwbar,
      qptr => accessQueueLength_qptr,
      wdata => accessQueueLength_wdata,
      rdata => accessQueueLength_rdata,
      start_req => accessQueueLength_start_req,
      start_ack => accessQueueLength_start_ack,
      fin_req => accessQueueLength_fin_req,
      fin_ack => accessQueueLength_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryWord_call_reqs => accessMemoryWord_call_reqs(2 downto 2),
      accessMemoryWord_call_acks => accessMemoryWord_call_acks(2 downto 2),
      accessMemoryWord_call_data => accessMemoryWord_call_data(506 downto 338),
      accessMemoryWord_call_tag => accessMemoryWord_call_tag(2 downto 2),
      accessMemoryWord_return_reqs => accessMemoryWord_return_reqs(2 downto 2),
      accessMemoryWord_return_acks => accessMemoryWord_return_acks(2 downto 2),
      accessMemoryWord_return_data => accessMemoryWord_return_data(95 downto 64),
      accessMemoryWord_return_tag => accessMemoryWord_return_tag(2 downto 2),
      tag_in => accessQueueLength_tag_in,
      tag_out => accessQueueLength_tag_out-- 
    ); -- 
  -- module accessQueueMisc
  accessQueueMisc_tag <= accessQueueMisc_in_args(104 downto 97);
  accessQueueMisc_rwbar <= accessQueueMisc_in_args(96 downto 96);
  accessQueueMisc_qptr <= accessQueueMisc_in_args(95 downto 32);
  accessQueueMisc_wdata <= accessQueueMisc_in_args(31 downto 0);
  accessQueueMisc_out_args <= accessQueueMisc_rdata ;
  -- call arbiter for module accessQueueMisc
  accessQueueMisc_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 105,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessQueueMisc_call_reqs,
      call_acks => accessQueueMisc_call_acks,
      return_reqs => accessQueueMisc_return_reqs,
      return_acks => accessQueueMisc_return_acks,
      call_data  => accessQueueMisc_call_data,
      call_tag  => accessQueueMisc_call_tag,
      return_tag  => accessQueueMisc_return_tag,
      call_mtag => accessQueueMisc_tag_in,
      return_mtag => accessQueueMisc_tag_out,
      return_data =>accessQueueMisc_return_data,
      call_mreq => accessQueueMisc_start_req,
      call_mack => accessQueueMisc_start_ack,
      return_mreq => accessQueueMisc_fin_req,
      return_mack => accessQueueMisc_fin_ack,
      call_mdata => accessQueueMisc_in_args,
      return_mdata => accessQueueMisc_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessQueueMisc_instance:accessQueueMisc-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => accessQueueMisc_tag,
      rwbar => accessQueueMisc_rwbar,
      qptr => accessQueueMisc_qptr,
      wdata => accessQueueMisc_wdata,
      rdata => accessQueueMisc_rdata,
      start_req => accessQueueMisc_start_req,
      start_ack => accessQueueMisc_start_ack,
      fin_req => accessQueueMisc_fin_req,
      fin_ack => accessQueueMisc_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryWord_call_reqs => accessMemoryWord_call_reqs(5 downto 5),
      accessMemoryWord_call_acks => accessMemoryWord_call_acks(5 downto 5),
      accessMemoryWord_call_data => accessMemoryWord_call_data(1013 downto 845),
      accessMemoryWord_call_tag => accessMemoryWord_call_tag(5 downto 5),
      accessMemoryWord_return_reqs => accessMemoryWord_return_reqs(5 downto 5),
      accessMemoryWord_return_acks => accessMemoryWord_return_acks(5 downto 5),
      accessMemoryWord_return_data => accessMemoryWord_return_data(191 downto 160),
      accessMemoryWord_return_tag => accessMemoryWord_return_tag(5 downto 5),
      tag_in => accessQueueMisc_tag_in,
      tag_out => accessQueueMisc_tag_out-- 
    ); -- 
  -- module accessQueueReadIndex
  accessQueueReadIndex_tag <= accessQueueReadIndex_in_args(104 downto 97);
  accessQueueReadIndex_rwbar <= accessQueueReadIndex_in_args(96 downto 96);
  accessQueueReadIndex_qptr <= accessQueueReadIndex_in_args(95 downto 32);
  accessQueueReadIndex_wdata <= accessQueueReadIndex_in_args(31 downto 0);
  accessQueueReadIndex_out_args <= accessQueueReadIndex_rdata ;
  -- call arbiter for module accessQueueReadIndex
  accessQueueReadIndex_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 105,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessQueueReadIndex_call_reqs,
      call_acks => accessQueueReadIndex_call_acks,
      return_reqs => accessQueueReadIndex_return_reqs,
      return_acks => accessQueueReadIndex_return_acks,
      call_data  => accessQueueReadIndex_call_data,
      call_tag  => accessQueueReadIndex_call_tag,
      return_tag  => accessQueueReadIndex_return_tag,
      call_mtag => accessQueueReadIndex_tag_in,
      return_mtag => accessQueueReadIndex_tag_out,
      return_data =>accessQueueReadIndex_return_data,
      call_mreq => accessQueueReadIndex_start_req,
      call_mack => accessQueueReadIndex_start_ack,
      return_mreq => accessQueueReadIndex_fin_req,
      return_mack => accessQueueReadIndex_fin_ack,
      call_mdata => accessQueueReadIndex_in_args,
      return_mdata => accessQueueReadIndex_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessQueueReadIndex_instance:accessQueueReadIndex-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => accessQueueReadIndex_tag,
      rwbar => accessQueueReadIndex_rwbar,
      qptr => accessQueueReadIndex_qptr,
      wdata => accessQueueReadIndex_wdata,
      rdata => accessQueueReadIndex_rdata,
      start_req => accessQueueReadIndex_start_req,
      start_ack => accessQueueReadIndex_start_ack,
      fin_req => accessQueueReadIndex_fin_req,
      fin_ack => accessQueueReadIndex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryWord_call_reqs => accessMemoryWord_call_reqs(4 downto 4),
      accessMemoryWord_call_acks => accessMemoryWord_call_acks(4 downto 4),
      accessMemoryWord_call_data => accessMemoryWord_call_data(844 downto 676),
      accessMemoryWord_call_tag => accessMemoryWord_call_tag(4 downto 4),
      accessMemoryWord_return_reqs => accessMemoryWord_return_reqs(4 downto 4),
      accessMemoryWord_return_acks => accessMemoryWord_return_acks(4 downto 4),
      accessMemoryWord_return_data => accessMemoryWord_return_data(159 downto 128),
      accessMemoryWord_return_tag => accessMemoryWord_return_tag(4 downto 4),
      tag_in => accessQueueReadIndex_tag_in,
      tag_out => accessQueueReadIndex_tag_out-- 
    ); -- 
  -- module accessQueueTotalMsgs
  accessQueueTotalMsgs_tag <= accessQueueTotalMsgs_in_args(104 downto 97);
  accessQueueTotalMsgs_rwbar <= accessQueueTotalMsgs_in_args(96 downto 96);
  accessQueueTotalMsgs_qptr <= accessQueueTotalMsgs_in_args(95 downto 32);
  accessQueueTotalMsgs_wdata <= accessQueueTotalMsgs_in_args(31 downto 0);
  accessQueueTotalMsgs_out_args <= accessQueueTotalMsgs_rdata ;
  -- call arbiter for module accessQueueTotalMsgs
  accessQueueTotalMsgs_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 105,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessQueueTotalMsgs_call_reqs,
      call_acks => accessQueueTotalMsgs_call_acks,
      return_reqs => accessQueueTotalMsgs_return_reqs,
      return_acks => accessQueueTotalMsgs_return_acks,
      call_data  => accessQueueTotalMsgs_call_data,
      call_tag  => accessQueueTotalMsgs_call_tag,
      return_tag  => accessQueueTotalMsgs_return_tag,
      call_mtag => accessQueueTotalMsgs_tag_in,
      return_mtag => accessQueueTotalMsgs_tag_out,
      return_data =>accessQueueTotalMsgs_return_data,
      call_mreq => accessQueueTotalMsgs_start_req,
      call_mack => accessQueueTotalMsgs_start_ack,
      return_mreq => accessQueueTotalMsgs_fin_req,
      return_mack => accessQueueTotalMsgs_fin_ack,
      call_mdata => accessQueueTotalMsgs_in_args,
      return_mdata => accessQueueTotalMsgs_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessQueueTotalMsgs_instance:accessQueueTotalMsgs-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => accessQueueTotalMsgs_tag,
      rwbar => accessQueueTotalMsgs_rwbar,
      qptr => accessQueueTotalMsgs_qptr,
      wdata => accessQueueTotalMsgs_wdata,
      rdata => accessQueueTotalMsgs_rdata,
      start_req => accessQueueTotalMsgs_start_req,
      start_ack => accessQueueTotalMsgs_start_ack,
      fin_req => accessQueueTotalMsgs_fin_req,
      fin_ack => accessQueueTotalMsgs_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryWord_call_reqs => accessMemoryWord_call_reqs(1 downto 1),
      accessMemoryWord_call_acks => accessMemoryWord_call_acks(1 downto 1),
      accessMemoryWord_call_data => accessMemoryWord_call_data(337 downto 169),
      accessMemoryWord_call_tag => accessMemoryWord_call_tag(1 downto 1),
      accessMemoryWord_return_reqs => accessMemoryWord_return_reqs(1 downto 1),
      accessMemoryWord_return_acks => accessMemoryWord_return_acks(1 downto 1),
      accessMemoryWord_return_data => accessMemoryWord_return_data(63 downto 32),
      accessMemoryWord_return_tag => accessMemoryWord_return_tag(1 downto 1),
      tag_in => accessQueueTotalMsgs_tag_in,
      tag_out => accessQueueTotalMsgs_tag_out-- 
    ); -- 
  -- module accessQueueWriteIndex
  accessQueueWriteIndex_tag <= accessQueueWriteIndex_in_args(104 downto 97);
  accessQueueWriteIndex_rwbar <= accessQueueWriteIndex_in_args(96 downto 96);
  accessQueueWriteIndex_qptr <= accessQueueWriteIndex_in_args(95 downto 32);
  accessQueueWriteIndex_wdata <= accessQueueWriteIndex_in_args(31 downto 0);
  accessQueueWriteIndex_out_args <= accessQueueWriteIndex_rdata ;
  -- call arbiter for module accessQueueWriteIndex
  accessQueueWriteIndex_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 105,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessQueueWriteIndex_call_reqs,
      call_acks => accessQueueWriteIndex_call_acks,
      return_reqs => accessQueueWriteIndex_return_reqs,
      return_acks => accessQueueWriteIndex_return_acks,
      call_data  => accessQueueWriteIndex_call_data,
      call_tag  => accessQueueWriteIndex_call_tag,
      return_tag  => accessQueueWriteIndex_return_tag,
      call_mtag => accessQueueWriteIndex_tag_in,
      return_mtag => accessQueueWriteIndex_tag_out,
      return_data =>accessQueueWriteIndex_return_data,
      call_mreq => accessQueueWriteIndex_start_req,
      call_mack => accessQueueWriteIndex_start_ack,
      return_mreq => accessQueueWriteIndex_fin_req,
      return_mack => accessQueueWriteIndex_fin_ack,
      call_mdata => accessQueueWriteIndex_in_args,
      return_mdata => accessQueueWriteIndex_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessQueueWriteIndex_instance:accessQueueWriteIndex-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => accessQueueWriteIndex_tag,
      rwbar => accessQueueWriteIndex_rwbar,
      qptr => accessQueueWriteIndex_qptr,
      wdata => accessQueueWriteIndex_wdata,
      rdata => accessQueueWriteIndex_rdata,
      start_req => accessQueueWriteIndex_start_req,
      start_ack => accessQueueWriteIndex_start_ack,
      fin_req => accessQueueWriteIndex_fin_req,
      fin_ack => accessQueueWriteIndex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryWord_call_reqs => accessMemoryWord_call_reqs(3 downto 3),
      accessMemoryWord_call_acks => accessMemoryWord_call_acks(3 downto 3),
      accessMemoryWord_call_data => accessMemoryWord_call_data(675 downto 507),
      accessMemoryWord_call_tag => accessMemoryWord_call_tag(3 downto 3),
      accessMemoryWord_return_reqs => accessMemoryWord_return_reqs(3 downto 3),
      accessMemoryWord_return_acks => accessMemoryWord_return_acks(3 downto 3),
      accessMemoryWord_return_data => accessMemoryWord_return_data(127 downto 96),
      accessMemoryWord_return_tag => accessMemoryWord_return_tag(3 downto 3),
      tag_in => accessQueueWriteIndex_tag_in,
      tag_out => accessQueueWriteIndex_tag_out-- 
    ); -- 
  -- module accessRegister
  accessRegister_rwbar <= accessRegister_in_args(44 downto 44);
  accessRegister_bmask <= accessRegister_in_args(43 downto 40);
  accessRegister_index <= accessRegister_in_args(39 downto 32);
  accessRegister_wdata <= accessRegister_in_args(31 downto 0);
  accessRegister_out_args <= accessRegister_rdata ;
  -- call arbiter for module accessRegister
  accessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 10,
      call_data_width => 45,
      return_data_width => 32,
      callee_tag_length => 4,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessRegister_call_reqs,
      call_acks => accessRegister_call_acks,
      return_reqs => accessRegister_return_reqs,
      return_acks => accessRegister_return_acks,
      call_data  => accessRegister_call_data,
      call_tag  => accessRegister_call_tag,
      return_tag  => accessRegister_return_tag,
      call_mtag => accessRegister_tag_in,
      return_mtag => accessRegister_tag_out,
      return_data =>accessRegister_return_data,
      call_mreq => accessRegister_start_req,
      call_mack => accessRegister_start_ack,
      return_mreq => accessRegister_fin_req,
      return_mack => accessRegister_fin_ack,
      call_mdata => accessRegister_in_args,
      return_mdata => accessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessRegister_instance:accessRegister-- 
    generic map(tag_length => 6)
    port map(-- 
      rwbar => accessRegister_rwbar,
      bmask => accessRegister_bmask,
      index => accessRegister_index,
      wdata => accessRegister_wdata,
      rdata => accessRegister_rdata,
      start_req => accessRegister_start_req,
      start_ack => accessRegister_start_ack,
      fin_req => accessRegister_fin_req,
      fin_ack => accessRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(7 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(7 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => accessRegister_tag_in,
      tag_out => accessRegister_tag_out-- 
    ); -- 
  -- module acquireLock
  acquireLock_tag <= acquireLock_in_args(71 downto 64);
  acquireLock_lock_address_pointer <= acquireLock_in_args(63 downto 0);
  acquireLock_out_args <= acquireLock_m_ok ;
  -- call arbiter for module acquireLock
  acquireLock_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 72,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireLock_call_reqs,
      call_acks => acquireLock_call_acks,
      return_reqs => acquireLock_return_reqs,
      return_acks => acquireLock_return_acks,
      call_data  => acquireLock_call_data,
      call_tag  => acquireLock_call_tag,
      return_tag  => acquireLock_return_tag,
      call_mtag => acquireLock_tag_in,
      return_mtag => acquireLock_tag_out,
      return_data =>acquireLock_return_data,
      call_mreq => acquireLock_start_req,
      call_mack => acquireLock_start_ack,
      return_mreq => acquireLock_fin_req,
      return_mack => acquireLock_fin_ack,
      call_mdata => acquireLock_in_args,
      return_mdata => acquireLock_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireLock_instance:acquireLock-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => acquireLock_tag,
      lock_address_pointer => acquireLock_lock_address_pointer,
      m_ok => acquireLock_m_ok,
      start_req => acquireLock_start_req,
      start_ack => acquireLock_start_ack,
      fin_req => acquireLock_fin_req,
      fin_ack => acquireLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryLdStub_call_reqs => accessMemoryLdStub_call_reqs(0 downto 0),
      accessMemoryLdStub_call_acks => accessMemoryLdStub_call_acks(0 downto 0),
      accessMemoryLdStub_call_data => accessMemoryLdStub_call_data(135 downto 0),
      accessMemoryLdStub_call_tag => accessMemoryLdStub_call_tag(0 downto 0),
      accessMemoryLdStub_return_reqs => accessMemoryLdStub_return_reqs(0 downto 0),
      accessMemoryLdStub_return_acks => accessMemoryLdStub_return_acks(0 downto 0),
      accessMemoryLdStub_return_data => accessMemoryLdStub_return_data(7 downto 0),
      accessMemoryLdStub_return_tag => accessMemoryLdStub_return_tag(0 downto 0),
      tag_in => acquireLock_tag_in,
      tag_out => acquireLock_tag_out-- 
    ); -- 
  -- module calculateAddress36
  calculateAddress36_addr_base <= calculateAddress36_in_args(127 downto 64);
  calculateAddress36_offset <= calculateAddress36_in_args(63 downto 0);
  calculateAddress36_out_args <= calculateAddress36_addr ;
  -- call arbiter for module calculateAddress36
  calculateAddress36_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 128,
      return_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => calculateAddress36_call_reqs,
      call_acks => calculateAddress36_call_acks,
      return_reqs => calculateAddress36_return_reqs,
      return_acks => calculateAddress36_return_acks,
      call_data  => calculateAddress36_call_data,
      call_tag  => calculateAddress36_call_tag,
      return_tag  => calculateAddress36_return_tag,
      call_mtag => calculateAddress36_tag_in,
      return_mtag => calculateAddress36_tag_out,
      return_data =>calculateAddress36_return_data,
      call_mreq => calculateAddress36_start_req,
      call_mack => calculateAddress36_start_ack,
      return_mreq => calculateAddress36_fin_req,
      return_mack => calculateAddress36_fin_ack,
      call_mdata => calculateAddress36_in_args,
      return_mdata => calculateAddress36_out_args,
      clk => clk, 
      reset => reset --
    ); --
  calculateAddress36_instance:calculateAddress36-- 
    generic map(tag_length => 3)
    port map(-- 
      addr_base => calculateAddress36_addr_base,
      offset => calculateAddress36_offset,
      addr => calculateAddress36_addr,
      start_req => calculateAddress36_start_req,
      start_ack => calculateAddress36_start_ack,
      fin_req => calculateAddress36_fin_req,
      fin_ack => calculateAddress36_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => calculateAddress36_tag_in,
      tag_out => calculateAddress36_tag_out-- 
    ); -- 
  -- module controlDaemon
  controlDaemon_instance:controlDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => controlDaemon_start_req,
      start_ack => controlDaemon_start_ack,
      fin_req => controlDaemon_fin_req,
      fin_ack => controlDaemon_fin_ack,
      clk => clk,
      reset => reset,
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      QUEUE_MONITOR_SIGNAL => QUEUE_MONITOR_SIGNAL,
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      NIC_INTR_pipe_write_req => NIC_INTR_pipe_write_req(0 downto 0),
      NIC_INTR_pipe_write_ack => NIC_INTR_pipe_write_ack(0 downto 0),
      NIC_INTR_pipe_write_data => NIC_INTR_pipe_write_data(0 downto 0),
      NIC_INTR_ENABLE_pipe_write_req => NIC_INTR_ENABLE_pipe_write_req(0 downto 0),
      NIC_INTR_ENABLE_pipe_write_ack => NIC_INTR_ENABLE_pipe_write_ack(0 downto 0),
      NIC_INTR_ENABLE_pipe_write_data => NIC_INTR_ENABLE_pipe_write_data(0 downto 0),
      MAC_ENABLE_pipe_write_req => MAC_ENABLE_pipe_write_req(0 downto 0),
      MAC_ENABLE_pipe_write_ack => MAC_ENABLE_pipe_write_ack(0 downto 0),
      MAC_ENABLE_pipe_write_data => MAC_ENABLE_pipe_write_data(0 downto 0),
      S_CONTROL_REGISTER_pipe_write_req => S_CONTROL_REGISTER_pipe_write_req(0 downto 0),
      S_CONTROL_REGISTER_pipe_write_ack => S_CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      S_CONTROL_REGISTER_pipe_write_data => S_CONTROL_REGISTER_pipe_write_data(31 downto 0),
      S_NUMBER_OF_SERVERS_pipe_write_req => S_NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      S_NUMBER_OF_SERVERS_pipe_write_ack => S_NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      S_NUMBER_OF_SERVERS_pipe_write_data => S_NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      NIC_INTR_INTERNAL_pipe_write_req => NIC_INTR_INTERNAL_pipe_write_req(0 downto 0),
      NIC_INTR_INTERNAL_pipe_write_ack => NIC_INTR_INTERNAL_pipe_write_ack(0 downto 0),
      NIC_INTR_INTERNAL_pipe_write_data => NIC_INTR_INTERNAL_pipe_write_data(0 downto 0),
      memory_access_lock_pipe_write_req => memory_access_lock_pipe_write_req(0 downto 0),
      memory_access_lock_pipe_write_ack => memory_access_lock_pipe_write_ack(0 downto 0),
      memory_access_lock_pipe_write_data => memory_access_lock_pipe_write_data(0 downto 0),
      accessRegister_call_reqs => accessRegister_call_reqs(3 downto 2),
      accessRegister_call_acks => accessRegister_call_acks(3 downto 2),
      accessRegister_call_data => accessRegister_call_data(179 downto 90),
      accessRegister_call_tag => accessRegister_call_tag(7 downto 4),
      accessRegister_return_reqs => accessRegister_return_reqs(3 downto 2),
      accessRegister_return_acks => accessRegister_return_acks(3 downto 2),
      accessRegister_return_data => accessRegister_return_data(127 downto 64),
      accessRegister_return_tag => accessRegister_return_tag(7 downto 4),
      setGlobalSignals_call_reqs => setGlobalSignals_call_reqs(0 downto 0),
      setGlobalSignals_call_acks => setGlobalSignals_call_acks(0 downto 0),
      setGlobalSignals_call_tag => setGlobalSignals_call_tag(0 downto 0),
      setGlobalSignals_return_reqs => setGlobalSignals_return_reqs(0 downto 0),
      setGlobalSignals_return_acks => setGlobalSignals_return_acks(0 downto 0),
      setGlobalSignals_return_tag => setGlobalSignals_return_tag(0 downto 0),
      tag_in => controlDaemon_tag_in,
      tag_out => controlDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  controlDaemon_tag_in <= (others => '0');
  controlDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => controlDaemon_start_req, start_ack => controlDaemon_start_ack,  fin_req => controlDaemon_fin_req,  fin_ack => controlDaemon_fin_ack);
  -- module doMemAccess
  doMemAccess_tag <= doMemAccess_in_args(202 downto 195);
  doMemAccess_opcode <= doMemAccess_in_args(194 downto 192);
  doMemAccess_base_addr <= doMemAccess_in_args(191 downto 128);
  doMemAccess_offset <= doMemAccess_in_args(127 downto 64);
  doMemAccess_wdata <= doMemAccess_in_args(63 downto 0);
  doMemAccess_out_args <= doMemAccess_rdata ;
  -- call arbiter for module doMemAccess
  doMemAccess_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 4,
      call_data_width => 203,
      return_data_width => 64,
      callee_tag_length => 3,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => doMemAccess_call_reqs,
      call_acks => doMemAccess_call_acks,
      return_reqs => doMemAccess_return_reqs,
      return_acks => doMemAccess_return_acks,
      call_data  => doMemAccess_call_data,
      call_tag  => doMemAccess_call_tag,
      return_tag  => doMemAccess_return_tag,
      call_mtag => doMemAccess_tag_in,
      return_mtag => doMemAccess_tag_out,
      return_data =>doMemAccess_return_data,
      call_mreq => doMemAccess_start_req,
      call_mack => doMemAccess_start_ack,
      return_mreq => doMemAccess_fin_req,
      return_mack => doMemAccess_fin_ack,
      call_mdata => doMemAccess_in_args,
      return_mdata => doMemAccess_out_args,
      clk => clk, 
      reset => reset --
    ); --
  doMemAccess_instance:doMemAccess-- 
    generic map(tag_length => 4)
    port map(-- 
      tag => doMemAccess_tag,
      opcode => doMemAccess_opcode,
      base_addr => doMemAccess_base_addr,
      offset => doMemAccess_offset,
      wdata => doMemAccess_wdata,
      rdata => doMemAccess_rdata,
      start_req => doMemAccess_start_req,
      start_ack => doMemAccess_start_ack,
      fin_req => doMemAccess_fin_req,
      fin_ack => doMemAccess_fin_ack,
      clk => clk,
      reset => reset,
      memory_access_lock_pipe_read_req => memory_access_lock_pipe_read_req(0 downto 0),
      memory_access_lock_pipe_read_ack => memory_access_lock_pipe_read_ack(0 downto 0),
      memory_access_lock_pipe_read_data => memory_access_lock_pipe_read_data(0 downto 0),
      memory_access_lock_pipe_write_req => memory_access_lock_pipe_write_req(1 downto 1),
      memory_access_lock_pipe_write_ack => memory_access_lock_pipe_write_ack(1 downto 1),
      memory_access_lock_pipe_write_data => memory_access_lock_pipe_write_data(1 downto 1),
      accessMemoryByteBase_call_reqs => accessMemoryByteBase_call_reqs(0 downto 0),
      accessMemoryByteBase_call_acks => accessMemoryByteBase_call_acks(0 downto 0),
      accessMemoryByteBase_call_data => accessMemoryByteBase_call_data(145 downto 0),
      accessMemoryByteBase_call_tag => accessMemoryByteBase_call_tag(1 downto 0),
      accessMemoryByteBase_return_reqs => accessMemoryByteBase_return_reqs(0 downto 0),
      accessMemoryByteBase_return_acks => accessMemoryByteBase_return_acks(0 downto 0),
      accessMemoryByteBase_return_data => accessMemoryByteBase_return_data(7 downto 0),
      accessMemoryByteBase_return_tag => accessMemoryByteBase_return_tag(1 downto 0),
      accessMemoryWordBase_call_reqs => accessMemoryWordBase_call_reqs(0 downto 0),
      accessMemoryWordBase_call_acks => accessMemoryWordBase_call_acks(0 downto 0),
      accessMemoryWordBase_call_data => accessMemoryWordBase_call_data(169 downto 0),
      accessMemoryWordBase_call_tag => accessMemoryWordBase_call_tag(0 downto 0),
      accessMemoryWordBase_return_reqs => accessMemoryWordBase_return_reqs(0 downto 0),
      accessMemoryWordBase_return_acks => accessMemoryWordBase_return_acks(0 downto 0),
      accessMemoryWordBase_return_data => accessMemoryWordBase_return_data(31 downto 0),
      accessMemoryWordBase_return_tag => accessMemoryWordBase_return_tag(0 downto 0),
      accessMemoryDwordBase_call_reqs => accessMemoryDwordBase_call_reqs(0 downto 0),
      accessMemoryDwordBase_call_acks => accessMemoryDwordBase_call_acks(0 downto 0),
      accessMemoryDwordBase_call_data => accessMemoryDwordBase_call_data(201 downto 0),
      accessMemoryDwordBase_call_tag => accessMemoryDwordBase_call_tag(0 downto 0),
      accessMemoryDwordBase_return_reqs => accessMemoryDwordBase_return_reqs(0 downto 0),
      accessMemoryDwordBase_return_acks => accessMemoryDwordBase_return_acks(0 downto 0),
      accessMemoryDwordBase_return_data => accessMemoryDwordBase_return_data(63 downto 0),
      accessMemoryDwordBase_return_tag => accessMemoryDwordBase_return_tag(0 downto 0),
      tag_in => doMemAccess_tag_in,
      tag_out => doMemAccess_tag_out-- 
    ); -- 
  -- module getQueueBufPointer
  getQueueBufPointer_queue_type <= getQueueBufPointer_in_args(9 downto 8);
  getQueueBufPointer_server_id <= getQueueBufPointer_in_args(7 downto 0);
  getQueueBufPointer_out_args <= getQueueBufPointer_qptr ;
  -- call arbiter for module getQueueBufPointer
  getQueueBufPointer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 10,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueBufPointer_call_reqs,
      call_acks => getQueueBufPointer_call_acks,
      return_reqs => getQueueBufPointer_return_reqs,
      return_acks => getQueueBufPointer_return_acks,
      call_data  => getQueueBufPointer_call_data,
      call_tag  => getQueueBufPointer_call_tag,
      return_tag  => getQueueBufPointer_return_tag,
      call_mtag => getQueueBufPointer_tag_in,
      return_mtag => getQueueBufPointer_tag_out,
      return_data =>getQueueBufPointer_return_data,
      call_mreq => getQueueBufPointer_start_req,
      call_mack => getQueueBufPointer_start_ack,
      return_mreq => getQueueBufPointer_fin_req,
      return_mack => getQueueBufPointer_fin_ack,
      call_mdata => getQueueBufPointer_in_args,
      return_mdata => getQueueBufPointer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueBufPointer_instance:getQueueBufPointer-- 
    generic map(tag_length => 3)
    port map(-- 
      queue_type => getQueueBufPointer_queue_type,
      server_id => getQueueBufPointer_server_id,
      qptr => getQueueBufPointer_qptr,
      start_req => getQueueBufPointer_start_req,
      start_ack => getQueueBufPointer_start_ack,
      fin_req => getQueueBufPointer_fin_req,
      fin_ack => getQueueBufPointer_fin_ack,
      clk => clk,
      reset => reset,
      accessRegister_call_reqs => accessRegister_call_reqs(7 downto 7),
      accessRegister_call_acks => accessRegister_call_acks(7 downto 7),
      accessRegister_call_data => accessRegister_call_data(359 downto 315),
      accessRegister_call_tag => accessRegister_call_tag(15 downto 14),
      accessRegister_return_reqs => accessRegister_return_reqs(7 downto 7),
      accessRegister_return_acks => accessRegister_return_acks(7 downto 7),
      accessRegister_return_data => accessRegister_return_data(255 downto 224),
      accessRegister_return_tag => accessRegister_return_tag(15 downto 14),
      tag_in => getQueueBufPointer_tag_in,
      tag_out => getQueueBufPointer_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_tag <= getQueueElement_in_args(103 downto 96);
  getQueueElement_buf_base_addr <= getQueueElement_in_args(95 downto 32);
  getQueueElement_read_index <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 104,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => getQueueElement_tag,
      buf_base_addr => getQueueElement_buf_base_addr,
      read_index => getQueueElement_read_index,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueElement_call_reqs => accessQueueElement_call_reqs(1 downto 1),
      accessQueueElement_call_acks => accessQueueElement_call_acks(1 downto 1),
      accessQueueElement_call_data => accessQueueElement_call_data(337 downto 169),
      accessQueueElement_call_tag => accessQueueElement_call_tag(1 downto 1),
      accessQueueElement_return_reqs => accessQueueElement_return_reqs(1 downto 1),
      accessQueueElement_return_acks => accessQueueElement_return_acks(1 downto 1),
      accessQueueElement_return_data => accessQueueElement_return_data(127 downto 64),
      accessQueueElement_return_tag => accessQueueElement_return_tag(1 downto 1),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueueLength
  getQueueLength_tag <= getQueueLength_in_args(71 downto 64);
  getQueueLength_q_base_address <= getQueueLength_in_args(63 downto 0);
  getQueueLength_out_args <= getQueueLength_queue_length ;
  -- call arbiter for module getQueueLength
  getQueueLength_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 72,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueLength_call_reqs,
      call_acks => getQueueLength_call_acks,
      return_reqs => getQueueLength_return_reqs,
      return_acks => getQueueLength_return_acks,
      call_data  => getQueueLength_call_data,
      call_tag  => getQueueLength_call_tag,
      return_tag  => getQueueLength_return_tag,
      call_mtag => getQueueLength_tag_in,
      return_mtag => getQueueLength_tag_out,
      return_data =>getQueueLength_return_data,
      call_mreq => getQueueLength_start_req,
      call_mack => getQueueLength_start_ack,
      return_mreq => getQueueLength_fin_req,
      return_mack => getQueueLength_fin_ack,
      call_mdata => getQueueLength_in_args,
      return_mdata => getQueueLength_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueLength_instance:getQueueLength-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => getQueueLength_tag,
      q_base_address => getQueueLength_q_base_address,
      queue_length => getQueueLength_queue_length,
      start_req => getQueueLength_start_req,
      start_ack => getQueueLength_start_ack,
      fin_req => getQueueLength_fin_req,
      fin_ack => getQueueLength_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueLength_call_reqs => accessQueueLength_call_reqs(0 downto 0),
      accessQueueLength_call_acks => accessQueueLength_call_acks(0 downto 0),
      accessQueueLength_call_data => accessQueueLength_call_data(104 downto 0),
      accessQueueLength_call_tag => accessQueueLength_call_tag(0 downto 0),
      accessQueueLength_return_reqs => accessQueueLength_return_reqs(0 downto 0),
      accessQueueLength_return_acks => accessQueueLength_return_acks(0 downto 0),
      accessQueueLength_return_data => accessQueueLength_return_data(31 downto 0),
      accessQueueLength_return_tag => accessQueueLength_return_tag(0 downto 0),
      tag_in => getQueueLength_tag_in,
      tag_out => getQueueLength_tag_out-- 
    ); -- 
  -- module getQueueLockPointer
  getQueueLockPointer_queue_type <= getQueueLockPointer_in_args(9 downto 8);
  getQueueLockPointer_server_id <= getQueueLockPointer_in_args(7 downto 0);
  getQueueLockPointer_out_args <= getQueueLockPointer_qptr ;
  -- call arbiter for module getQueueLockPointer
  getQueueLockPointer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 10,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueLockPointer_call_reqs,
      call_acks => getQueueLockPointer_call_acks,
      return_reqs => getQueueLockPointer_return_reqs,
      return_acks => getQueueLockPointer_return_acks,
      call_data  => getQueueLockPointer_call_data,
      call_tag  => getQueueLockPointer_call_tag,
      return_tag  => getQueueLockPointer_return_tag,
      call_mtag => getQueueLockPointer_tag_in,
      return_mtag => getQueueLockPointer_tag_out,
      return_data =>getQueueLockPointer_return_data,
      call_mreq => getQueueLockPointer_start_req,
      call_mack => getQueueLockPointer_start_ack,
      return_mreq => getQueueLockPointer_fin_req,
      return_mack => getQueueLockPointer_fin_ack,
      call_mdata => getQueueLockPointer_in_args,
      return_mdata => getQueueLockPointer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueLockPointer_instance:getQueueLockPointer-- 
    generic map(tag_length => 3)
    port map(-- 
      queue_type => getQueueLockPointer_queue_type,
      server_id => getQueueLockPointer_server_id,
      qptr => getQueueLockPointer_qptr,
      start_req => getQueueLockPointer_start_req,
      start_ack => getQueueLockPointer_start_ack,
      fin_req => getQueueLockPointer_fin_req,
      fin_ack => getQueueLockPointer_fin_ack,
      clk => clk,
      reset => reset,
      accessRegister_call_reqs => accessRegister_call_reqs(8 downto 8),
      accessRegister_call_acks => accessRegister_call_acks(8 downto 8),
      accessRegister_call_data => accessRegister_call_data(404 downto 360),
      accessRegister_call_tag => accessRegister_call_tag(17 downto 16),
      accessRegister_return_reqs => accessRegister_return_reqs(8 downto 8),
      accessRegister_return_acks => accessRegister_return_acks(8 downto 8),
      accessRegister_return_data => accessRegister_return_data(287 downto 256),
      accessRegister_return_tag => accessRegister_return_tag(17 downto 16),
      tag_in => getQueueLockPointer_tag_in,
      tag_out => getQueueLockPointer_tag_out-- 
    ); -- 
  -- module getQueuePointer
  getQueuePointer_queue_type <= getQueuePointer_in_args(9 downto 8);
  getQueuePointer_server_id <= getQueuePointer_in_args(7 downto 0);
  getQueuePointer_out_args <= getQueuePointer_qptr ;
  -- call arbiter for module getQueuePointer
  getQueuePointer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 10,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointer_call_reqs,
      call_acks => getQueuePointer_call_acks,
      return_reqs => getQueuePointer_return_reqs,
      return_acks => getQueuePointer_return_acks,
      call_data  => getQueuePointer_call_data,
      call_tag  => getQueuePointer_call_tag,
      return_tag  => getQueuePointer_return_tag,
      call_mtag => getQueuePointer_tag_in,
      return_mtag => getQueuePointer_tag_out,
      return_data =>getQueuePointer_return_data,
      call_mreq => getQueuePointer_start_req,
      call_mack => getQueuePointer_start_ack,
      return_mreq => getQueuePointer_fin_req,
      return_mack => getQueuePointer_fin_ack,
      call_mdata => getQueuePointer_in_args,
      return_mdata => getQueuePointer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointer_instance:getQueuePointer-- 
    generic map(tag_length => 3)
    port map(-- 
      queue_type => getQueuePointer_queue_type,
      server_id => getQueuePointer_server_id,
      qptr => getQueuePointer_qptr,
      start_req => getQueuePointer_start_req,
      start_ack => getQueuePointer_start_ack,
      fin_req => getQueuePointer_fin_req,
      fin_ack => getQueuePointer_fin_ack,
      clk => clk,
      reset => reset,
      accessRegister_call_reqs => accessRegister_call_reqs(9 downto 9),
      accessRegister_call_acks => accessRegister_call_acks(9 downto 9),
      accessRegister_call_data => accessRegister_call_data(449 downto 405),
      accessRegister_call_tag => accessRegister_call_tag(19 downto 18),
      accessRegister_return_reqs => accessRegister_return_reqs(9 downto 9),
      accessRegister_return_acks => accessRegister_return_acks(9 downto 9),
      accessRegister_return_data => accessRegister_return_data(319 downto 288),
      accessRegister_return_tag => accessRegister_return_tag(19 downto 18),
      tag_in => getQueuePointer_tag_in,
      tag_out => getQueuePointer_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_tag <= getQueuePointers_in_args(71 downto 64);
  getQueuePointers_q_base_address <= getQueuePointers_in_args(63 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 72,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => getQueuePointers_tag,
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueReadIndex_call_reqs => accessQueueReadIndex_call_reqs(0 downto 0),
      accessQueueReadIndex_call_acks => accessQueueReadIndex_call_acks(0 downto 0),
      accessQueueReadIndex_call_data => accessQueueReadIndex_call_data(104 downto 0),
      accessQueueReadIndex_call_tag => accessQueueReadIndex_call_tag(0 downto 0),
      accessQueueReadIndex_return_reqs => accessQueueReadIndex_return_reqs(0 downto 0),
      accessQueueReadIndex_return_acks => accessQueueReadIndex_return_acks(0 downto 0),
      accessQueueReadIndex_return_data => accessQueueReadIndex_return_data(31 downto 0),
      accessQueueReadIndex_return_tag => accessQueueReadIndex_return_tag(0 downto 0),
      accessQueueWriteIndex_call_reqs => accessQueueWriteIndex_call_reqs(0 downto 0),
      accessQueueWriteIndex_call_acks => accessQueueWriteIndex_call_acks(0 downto 0),
      accessQueueWriteIndex_call_data => accessQueueWriteIndex_call_data(104 downto 0),
      accessQueueWriteIndex_call_tag => accessQueueWriteIndex_call_tag(0 downto 0),
      accessQueueWriteIndex_return_reqs => accessQueueWriteIndex_return_reqs(0 downto 0),
      accessQueueWriteIndex_return_acks => accessQueueWriteIndex_return_acks(0 downto 0),
      accessQueueWriteIndex_return_data => accessQueueWriteIndex_return_data(31 downto 0),
      accessQueueWriteIndex_return_tag => accessQueueWriteIndex_return_tag(0 downto 0),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTotalMessages
  getTotalMessages_tag <= getTotalMessages_in_args(71 downto 64);
  getTotalMessages_q_base_address <= getTotalMessages_in_args(63 downto 0);
  getTotalMessages_out_args <= getTotalMessages_total_msgs ;
  -- call arbiter for module getTotalMessages
  getTotalMessages_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 72,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTotalMessages_call_reqs,
      call_acks => getTotalMessages_call_acks,
      return_reqs => getTotalMessages_return_reqs,
      return_acks => getTotalMessages_return_acks,
      call_data  => getTotalMessages_call_data,
      call_tag  => getTotalMessages_call_tag,
      return_tag  => getTotalMessages_return_tag,
      call_mtag => getTotalMessages_tag_in,
      return_mtag => getTotalMessages_tag_out,
      return_data =>getTotalMessages_return_data,
      call_mreq => getTotalMessages_start_req,
      call_mack => getTotalMessages_start_ack,
      return_mreq => getTotalMessages_fin_req,
      return_mack => getTotalMessages_fin_ack,
      call_mdata => getTotalMessages_in_args,
      return_mdata => getTotalMessages_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTotalMessages_instance:getTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => getTotalMessages_tag,
      q_base_address => getTotalMessages_q_base_address,
      total_msgs => getTotalMessages_total_msgs,
      start_req => getTotalMessages_start_req,
      start_ack => getTotalMessages_start_ack,
      fin_req => getTotalMessages_fin_req,
      fin_ack => getTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueTotalMsgs_call_reqs => accessQueueTotalMsgs_call_reqs(0 downto 0),
      accessQueueTotalMsgs_call_acks => accessQueueTotalMsgs_call_acks(0 downto 0),
      accessQueueTotalMsgs_call_data => accessQueueTotalMsgs_call_data(104 downto 0),
      accessQueueTotalMsgs_call_tag => accessQueueTotalMsgs_call_tag(0 downto 0),
      accessQueueTotalMsgs_return_reqs => accessQueueTotalMsgs_return_reqs(0 downto 0),
      accessQueueTotalMsgs_return_acks => accessQueueTotalMsgs_return_acks(0 downto 0),
      accessQueueTotalMsgs_return_data => accessQueueTotalMsgs_return_data(31 downto 0),
      accessQueueTotalMsgs_return_tag => accessQueueTotalMsgs_return_tag(0 downto 0),
      tag_in => getTotalMessages_tag_in,
      tag_out => getTotalMessages_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_tag <= getTxPacketPointerFromServer_in_args(15 downto 8);
  getTxPacketPointerFromServer_server_index <= getTxPacketPointerFromServer_in_args(7 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 16,
      return_data_width => 65,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => getTxPacketPointerFromServer_tag,
      server_index => getTxPacketPointerFromServer_server_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(17 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(64 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module incrementNumberOfPacketsReceived
  -- call arbiter for module incrementNumberOfPacketsReceived
  incrementNumberOfPacketsReceived_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => incrementNumberOfPacketsReceived_call_reqs,
      call_acks => incrementNumberOfPacketsReceived_call_acks,
      return_reqs => incrementNumberOfPacketsReceived_return_reqs,
      return_acks => incrementNumberOfPacketsReceived_return_acks,
      call_tag  => incrementNumberOfPacketsReceived_call_tag,
      return_tag  => incrementNumberOfPacketsReceived_return_tag,
      call_mtag => incrementNumberOfPacketsReceived_tag_in,
      return_mtag => incrementNumberOfPacketsReceived_tag_out,
      call_mreq => incrementNumberOfPacketsReceived_start_req,
      call_mack => incrementNumberOfPacketsReceived_start_ack,
      return_mreq => incrementNumberOfPacketsReceived_fin_req,
      return_mack => incrementNumberOfPacketsReceived_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  incrementNumberOfPacketsReceived_instance:incrementNumberOfPacketsReceived-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => incrementNumberOfPacketsReceived_start_req,
      start_ack => incrementNumberOfPacketsReceived_start_ack,
      fin_req => incrementNumberOfPacketsReceived_fin_req,
      fin_ack => incrementNumberOfPacketsReceived_fin_ack,
      clk => clk,
      reset => reset,
      incrementRegister_call_reqs => incrementRegister_call_reqs(1 downto 1),
      incrementRegister_call_acks => incrementRegister_call_acks(1 downto 1),
      incrementRegister_call_data => incrementRegister_call_data(15 downto 8),
      incrementRegister_call_tag => incrementRegister_call_tag(1 downto 1),
      incrementRegister_return_reqs => incrementRegister_return_reqs(1 downto 1),
      incrementRegister_return_acks => incrementRegister_return_acks(1 downto 1),
      incrementRegister_return_data => incrementRegister_return_data(63 downto 32),
      incrementRegister_return_tag => incrementRegister_return_tag(1 downto 1),
      tag_in => incrementNumberOfPacketsReceived_tag_in,
      tag_out => incrementNumberOfPacketsReceived_tag_out-- 
    ); -- 
  -- module incrementNumberOfPacketsTransmitted
  -- call arbiter for module incrementNumberOfPacketsTransmitted
  incrementNumberOfPacketsTransmitted_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => incrementNumberOfPacketsTransmitted_call_reqs,
      call_acks => incrementNumberOfPacketsTransmitted_call_acks,
      return_reqs => incrementNumberOfPacketsTransmitted_return_reqs,
      return_acks => incrementNumberOfPacketsTransmitted_return_acks,
      call_tag  => incrementNumberOfPacketsTransmitted_call_tag,
      return_tag  => incrementNumberOfPacketsTransmitted_return_tag,
      call_mtag => incrementNumberOfPacketsTransmitted_tag_in,
      return_mtag => incrementNumberOfPacketsTransmitted_tag_out,
      call_mreq => incrementNumberOfPacketsTransmitted_start_req,
      call_mack => incrementNumberOfPacketsTransmitted_start_ack,
      return_mreq => incrementNumberOfPacketsTransmitted_fin_req,
      return_mack => incrementNumberOfPacketsTransmitted_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  incrementNumberOfPacketsTransmitted_instance:incrementNumberOfPacketsTransmitted-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => incrementNumberOfPacketsTransmitted_start_req,
      start_ack => incrementNumberOfPacketsTransmitted_start_ack,
      fin_req => incrementNumberOfPacketsTransmitted_fin_req,
      fin_ack => incrementNumberOfPacketsTransmitted_fin_ack,
      clk => clk,
      reset => reset,
      incrementRegister_call_reqs => incrementRegister_call_reqs(0 downto 0),
      incrementRegister_call_acks => incrementRegister_call_acks(0 downto 0),
      incrementRegister_call_data => incrementRegister_call_data(7 downto 0),
      incrementRegister_call_tag => incrementRegister_call_tag(0 downto 0),
      incrementRegister_return_reqs => incrementRegister_return_reqs(0 downto 0),
      incrementRegister_return_acks => incrementRegister_return_acks(0 downto 0),
      incrementRegister_return_data => incrementRegister_return_data(31 downto 0),
      incrementRegister_return_tag => incrementRegister_return_tag(0 downto 0),
      tag_in => incrementNumberOfPacketsTransmitted_tag_in,
      tag_out => incrementNumberOfPacketsTransmitted_tag_out-- 
    ); -- 
  -- module incrementRegister
  incrementRegister_reg_index <= incrementRegister_in_args(7 downto 0);
  incrementRegister_out_args <= incrementRegister_incremented_value ;
  -- call arbiter for module incrementRegister
  incrementRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 8,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => incrementRegister_call_reqs,
      call_acks => incrementRegister_call_acks,
      return_reqs => incrementRegister_return_reqs,
      return_acks => incrementRegister_return_acks,
      call_data  => incrementRegister_call_data,
      call_tag  => incrementRegister_call_tag,
      return_tag  => incrementRegister_return_tag,
      call_mtag => incrementRegister_tag_in,
      return_mtag => incrementRegister_tag_out,
      return_data =>incrementRegister_return_data,
      call_mreq => incrementRegister_start_req,
      call_mack => incrementRegister_start_ack,
      return_mreq => incrementRegister_fin_req,
      return_mack => incrementRegister_fin_ack,
      call_mdata => incrementRegister_in_args,
      return_mdata => incrementRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  incrementRegister_instance:incrementRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      reg_index => incrementRegister_reg_index,
      incremented_value => incrementRegister_incremented_value,
      start_req => incrementRegister_start_req,
      start_ack => incrementRegister_start_ack,
      fin_req => incrementRegister_fin_req,
      fin_ack => incrementRegister_fin_ack,
      clk => clk,
      reset => reset,
      accessRegister_call_reqs => accessRegister_call_reqs(6 downto 6),
      accessRegister_call_acks => accessRegister_call_acks(6 downto 6),
      accessRegister_call_data => accessRegister_call_data(314 downto 270),
      accessRegister_call_tag => accessRegister_call_tag(13 downto 12),
      accessRegister_return_reqs => accessRegister_return_reqs(6 downto 6),
      accessRegister_return_acks => accessRegister_return_acks(6 downto 6),
      accessRegister_return_data => accessRegister_return_data(223 downto 192),
      accessRegister_return_tag => accessRegister_return_tag(13 downto 12),
      tag_in => incrementRegister_tag_in,
      tag_out => incrementRegister_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_tag <= loadBuffer_in_args(87 downto 80);
  loadBuffer_max_addr_offset <= loadBuffer_in_args(79 downto 64);
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(63 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 88,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => loadBuffer_tag,
      max_addr_offset => loadBuffer_max_addr_offset,
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(71 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(15 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(103 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(19 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(106 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      S_CONTROL_REGISTER => S_CONTROL_REGISTER,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      accessRegister_call_reqs => accessRegister_call_reqs(1 downto 0),
      accessRegister_call_acks => accessRegister_call_acks(1 downto 0),
      accessRegister_call_data => accessRegister_call_data(89 downto 0),
      accessRegister_call_tag => accessRegister_call_tag(3 downto 0),
      accessRegister_return_reqs => accessRegister_return_reqs(1 downto 0),
      accessRegister_return_acks => accessRegister_return_acks(1 downto 0),
      accessRegister_return_data => accessRegister_return_data(63 downto 0),
      accessRegister_return_tag => accessRegister_return_tag(3 downto 0),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module popFromQueue
  popFromQueue_tag <= popFromQueue_in_args(17 downto 10);
  popFromQueue_queue_type <= popFromQueue_in_args(9 downto 8);
  popFromQueue_server_id <= popFromQueue_in_args(7 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 18,
      return_data_width => 65,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => popFromQueue_tag,
      queue_type => popFromQueue_queue_type,
      server_id => popFromQueue_server_id,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      QUEUE_MONITOR_SIGNAL_pipe_write_req => QUEUE_MONITOR_SIGNAL_pipe_write_req(1 downto 1),
      QUEUE_MONITOR_SIGNAL_pipe_write_ack => QUEUE_MONITOR_SIGNAL_pipe_write_ack(1 downto 1),
      QUEUE_MONITOR_SIGNAL_pipe_write_data => QUEUE_MONITOR_SIGNAL_pipe_write_data(63 downto 32),
      getQueuePointer_call_reqs => getQueuePointer_call_reqs(1 downto 1),
      getQueuePointer_call_acks => getQueuePointer_call_acks(1 downto 1),
      getQueuePointer_call_data => getQueuePointer_call_data(19 downto 10),
      getQueuePointer_call_tag => getQueuePointer_call_tag(1 downto 1),
      getQueuePointer_return_reqs => getQueuePointer_return_reqs(1 downto 1),
      getQueuePointer_return_acks => getQueuePointer_return_acks(1 downto 1),
      getQueuePointer_return_data => getQueuePointer_return_data(127 downto 64),
      getQueuePointer_return_tag => getQueuePointer_return_tag(1 downto 1),
      accessQueueMisc_call_reqs => accessQueueMisc_call_reqs(0 downto 0),
      accessQueueMisc_call_acks => accessQueueMisc_call_acks(0 downto 0),
      accessQueueMisc_call_data => accessQueueMisc_call_data(104 downto 0),
      accessQueueMisc_call_tag => accessQueueMisc_call_tag(0 downto 0),
      accessQueueMisc_return_reqs => accessQueueMisc_return_reqs(0 downto 0),
      accessQueueMisc_return_acks => accessQueueMisc_return_acks(0 downto 0),
      accessQueueMisc_return_data => accessQueueMisc_return_data(31 downto 0),
      accessQueueMisc_return_tag => accessQueueMisc_return_tag(0 downto 0),
      getQueueLockPointer_call_reqs => getQueueLockPointer_call_reqs(1 downto 1),
      getQueueLockPointer_call_acks => getQueueLockPointer_call_acks(1 downto 1),
      getQueueLockPointer_call_data => getQueueLockPointer_call_data(19 downto 10),
      getQueueLockPointer_call_tag => getQueueLockPointer_call_tag(1 downto 1),
      getQueueLockPointer_return_reqs => getQueueLockPointer_return_reqs(1 downto 1),
      getQueueLockPointer_return_acks => getQueueLockPointer_return_acks(1 downto 1),
      getQueueLockPointer_return_data => getQueueLockPointer_return_data(127 downto 64),
      getQueueLockPointer_return_tag => getQueueLockPointer_return_tag(1 downto 1),
      acquireLock_call_reqs => acquireLock_call_reqs(1 downto 1),
      acquireLock_call_acks => acquireLock_call_acks(1 downto 1),
      acquireLock_call_data => acquireLock_call_data(143 downto 72),
      acquireLock_call_tag => acquireLock_call_tag(1 downto 1),
      acquireLock_return_reqs => acquireLock_return_reqs(1 downto 1),
      acquireLock_return_acks => acquireLock_return_acks(1 downto 1),
      acquireLock_return_data => acquireLock_return_data(1 downto 1),
      acquireLock_return_tag => acquireLock_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(143 downto 72),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      getQueueLength_call_reqs => getQueueLength_call_reqs(1 downto 1),
      getQueueLength_call_acks => getQueueLength_call_acks(1 downto 1),
      getQueueLength_call_data => getQueueLength_call_data(143 downto 72),
      getQueueLength_call_tag => getQueueLength_call_tag(1 downto 1),
      getQueueLength_return_reqs => getQueueLength_return_reqs(1 downto 1),
      getQueueLength_return_acks => getQueueLength_return_acks(1 downto 1),
      getQueueLength_return_data => getQueueLength_return_data(63 downto 32),
      getQueueLength_return_tag => getQueueLength_return_tag(1 downto 1),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(1 downto 1),
      getTotalMessages_call_acks => getTotalMessages_call_acks(1 downto 1),
      getTotalMessages_call_data => getTotalMessages_call_data(143 downto 72),
      getTotalMessages_call_tag => getTotalMessages_call_tag(1 downto 1),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(1 downto 1),
      getTotalMessages_return_acks => getTotalMessages_return_acks(1 downto 1),
      getTotalMessages_return_data => getTotalMessages_return_data(63 downto 32),
      getTotalMessages_return_tag => getTotalMessages_return_tag(1 downto 1),
      getQueueBufPointer_call_reqs => getQueueBufPointer_call_reqs(1 downto 1),
      getQueueBufPointer_call_acks => getQueueBufPointer_call_acks(1 downto 1),
      getQueueBufPointer_call_data => getQueueBufPointer_call_data(19 downto 10),
      getQueueBufPointer_call_tag => getQueueBufPointer_call_tag(1 downto 1),
      getQueueBufPointer_return_reqs => getQueueBufPointer_return_reqs(1 downto 1),
      getQueueBufPointer_return_acks => getQueueBufPointer_return_acks(1 downto 1),
      getQueueBufPointer_return_data => getQueueBufPointer_return_data(127 downto 64),
      getQueueBufPointer_return_tag => getQueueBufPointer_return_tag(1 downto 1),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(103 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(63 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(271 downto 136),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      setTotalMessages_call_reqs => setTotalMessages_call_reqs(1 downto 1),
      setTotalMessages_call_acks => setTotalMessages_call_acks(1 downto 1),
      setTotalMessages_call_data => setTotalMessages_call_data(207 downto 104),
      setTotalMessages_call_tag => setTotalMessages_call_tag(1 downto 1),
      setTotalMessages_return_reqs => setTotalMessages_return_reqs(1 downto 1),
      setTotalMessages_return_acks => setTotalMessages_return_acks(1 downto 1),
      setTotalMessages_return_tag => setTotalMessages_return_tag(1 downto 1),
      releaseLock_call_reqs => releaseLock_call_reqs(1 downto 1),
      releaseLock_call_acks => releaseLock_call_acks(1 downto 1),
      releaseLock_call_data => releaseLock_call_data(143 downto 72),
      releaseLock_call_tag => releaseLock_call_tag(1 downto 1),
      releaseLock_return_reqs => releaseLock_return_reqs(1 downto 1),
      releaseLock_return_acks => releaseLock_return_acks(1 downto 1),
      releaseLock_return_tag => releaseLock_return_tag(1 downto 1),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_tag <= populateRxQueue_in_args(71 downto 64);
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(63 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 72,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => populateRxQueue_tag,
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      S_NUMBER_OF_SERVERS => S_NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(15 downto 8),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(245 downto 164),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      incrementNumberOfPacketsReceived_call_reqs => incrementNumberOfPacketsReceived_call_reqs(0 downto 0),
      incrementNumberOfPacketsReceived_call_acks => incrementNumberOfPacketsReceived_call_acks(0 downto 0),
      incrementNumberOfPacketsReceived_call_tag => incrementNumberOfPacketsReceived_call_tag(0 downto 0),
      incrementNumberOfPacketsReceived_return_reqs => incrementNumberOfPacketsReceived_return_reqs(0 downto 0),
      incrementNumberOfPacketsReceived_return_acks => incrementNumberOfPacketsReceived_return_acks(0 downto 0),
      incrementNumberOfPacketsReceived_return_tag => incrementNumberOfPacketsReceived_return_tag(0 downto 0),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module pushIntoQueue
  pushIntoQueue_tag <= pushIntoQueue_in_args(81 downto 74);
  pushIntoQueue_queue_type <= pushIntoQueue_in_args(73 downto 72);
  pushIntoQueue_server_id <= pushIntoQueue_in_args(71 downto 64);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(63 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 82,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => pushIntoQueue_tag,
      queue_type => pushIntoQueue_queue_type,
      server_id => pushIntoQueue_server_id,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      QUEUE_MONITOR_SIGNAL_pipe_write_req => QUEUE_MONITOR_SIGNAL_pipe_write_req(0 downto 0),
      QUEUE_MONITOR_SIGNAL_pipe_write_ack => QUEUE_MONITOR_SIGNAL_pipe_write_ack(0 downto 0),
      QUEUE_MONITOR_SIGNAL_pipe_write_data => QUEUE_MONITOR_SIGNAL_pipe_write_data(31 downto 0),
      getQueuePointer_call_reqs => getQueuePointer_call_reqs(0 downto 0),
      getQueuePointer_call_acks => getQueuePointer_call_acks(0 downto 0),
      getQueuePointer_call_data => getQueuePointer_call_data(9 downto 0),
      getQueuePointer_call_tag => getQueuePointer_call_tag(0 downto 0),
      getQueuePointer_return_reqs => getQueuePointer_return_reqs(0 downto 0),
      getQueuePointer_return_acks => getQueuePointer_return_acks(0 downto 0),
      getQueuePointer_return_data => getQueuePointer_return_data(63 downto 0),
      getQueuePointer_return_tag => getQueuePointer_return_tag(0 downto 0),
      accessMemoryWord_call_reqs => accessMemoryWord_call_reqs(0 downto 0),
      accessMemoryWord_call_acks => accessMemoryWord_call_acks(0 downto 0),
      accessMemoryWord_call_data => accessMemoryWord_call_data(168 downto 0),
      accessMemoryWord_call_tag => accessMemoryWord_call_tag(0 downto 0),
      accessMemoryWord_return_reqs => accessMemoryWord_return_reqs(0 downto 0),
      accessMemoryWord_return_acks => accessMemoryWord_return_acks(0 downto 0),
      accessMemoryWord_return_data => accessMemoryWord_return_data(31 downto 0),
      accessMemoryWord_return_tag => accessMemoryWord_return_tag(0 downto 0),
      getQueueLockPointer_call_reqs => getQueueLockPointer_call_reqs(0 downto 0),
      getQueueLockPointer_call_acks => getQueueLockPointer_call_acks(0 downto 0),
      getQueueLockPointer_call_data => getQueueLockPointer_call_data(9 downto 0),
      getQueueLockPointer_call_tag => getQueueLockPointer_call_tag(0 downto 0),
      getQueueLockPointer_return_reqs => getQueueLockPointer_return_reqs(0 downto 0),
      getQueueLockPointer_return_acks => getQueueLockPointer_return_acks(0 downto 0),
      getQueueLockPointer_return_data => getQueueLockPointer_return_data(63 downto 0),
      getQueueLockPointer_return_tag => getQueueLockPointer_return_tag(0 downto 0),
      acquireLock_call_reqs => acquireLock_call_reqs(0 downto 0),
      acquireLock_call_acks => acquireLock_call_acks(0 downto 0),
      acquireLock_call_data => acquireLock_call_data(71 downto 0),
      acquireLock_call_tag => acquireLock_call_tag(0 downto 0),
      acquireLock_return_reqs => acquireLock_return_reqs(0 downto 0),
      acquireLock_return_acks => acquireLock_return_acks(0 downto 0),
      acquireLock_return_data => acquireLock_return_data(0 downto 0),
      acquireLock_return_tag => acquireLock_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      getQueueLength_call_reqs => getQueueLength_call_reqs(0 downto 0),
      getQueueLength_call_acks => getQueueLength_call_acks(0 downto 0),
      getQueueLength_call_data => getQueueLength_call_data(71 downto 0),
      getQueueLength_call_tag => getQueueLength_call_tag(0 downto 0),
      getQueueLength_return_reqs => getQueueLength_return_reqs(0 downto 0),
      getQueueLength_return_acks => getQueueLength_return_acks(0 downto 0),
      getQueueLength_return_data => getQueueLength_return_data(31 downto 0),
      getQueueLength_return_tag => getQueueLength_return_tag(0 downto 0),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(0 downto 0),
      getTotalMessages_call_acks => getTotalMessages_call_acks(0 downto 0),
      getTotalMessages_call_data => getTotalMessages_call_data(71 downto 0),
      getTotalMessages_call_tag => getTotalMessages_call_tag(0 downto 0),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(0 downto 0),
      getTotalMessages_return_acks => getTotalMessages_return_acks(0 downto 0),
      getTotalMessages_return_data => getTotalMessages_return_data(31 downto 0),
      getTotalMessages_return_tag => getTotalMessages_return_tag(0 downto 0),
      getQueueBufPointer_call_reqs => getQueueBufPointer_call_reqs(0 downto 0),
      getQueueBufPointer_call_acks => getQueueBufPointer_call_acks(0 downto 0),
      getQueueBufPointer_call_data => getQueueBufPointer_call_data(9 downto 0),
      getQueueBufPointer_call_tag => getQueueBufPointer_call_tag(0 downto 0),
      getQueueBufPointer_return_reqs => getQueueBufPointer_return_reqs(0 downto 0),
      getQueueBufPointer_return_acks => getQueueBufPointer_return_acks(0 downto 0),
      getQueueBufPointer_return_data => getQueueBufPointer_return_data(63 downto 0),
      getQueueBufPointer_return_tag => getQueueBufPointer_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(135 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      setTotalMessages_call_reqs => setTotalMessages_call_reqs(0 downto 0),
      setTotalMessages_call_acks => setTotalMessages_call_acks(0 downto 0),
      setTotalMessages_call_data => setTotalMessages_call_data(103 downto 0),
      setTotalMessages_call_tag => setTotalMessages_call_tag(0 downto 0),
      setTotalMessages_return_reqs => setTotalMessages_return_reqs(0 downto 0),
      setTotalMessages_return_acks => setTotalMessages_return_acks(0 downto 0),
      setTotalMessages_return_tag => setTotalMessages_return_tag(0 downto 0),
      releaseLock_call_reqs => releaseLock_call_reqs(0 downto 0),
      releaseLock_call_acks => releaseLock_call_acks(0 downto 0),
      releaseLock_call_data => releaseLock_call_data(71 downto 0),
      releaseLock_call_tag => releaseLock_call_tag(0 downto 0),
      releaseLock_return_reqs => releaseLock_return_reqs(0 downto 0),
      releaseLock_return_acks => releaseLock_return_acks(0 downto 0),
      releaseLock_return_tag => releaseLock_return_tag(0 downto 0),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(167 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseLock
  releaseLock_tag <= releaseLock_in_args(71 downto 64);
  releaseLock_lock_address_pointer <= releaseLock_in_args(63 downto 0);
  -- call arbiter for module releaseLock
  releaseLock_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 72,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseLock_call_reqs,
      call_acks => releaseLock_call_acks,
      return_reqs => releaseLock_return_reqs,
      return_acks => releaseLock_return_acks,
      call_data  => releaseLock_call_data,
      call_tag  => releaseLock_call_tag,
      return_tag  => releaseLock_return_tag,
      call_mtag => releaseLock_tag_in,
      return_mtag => releaseLock_tag_out,
      call_mreq => releaseLock_start_req,
      call_mack => releaseLock_start_ack,
      return_mreq => releaseLock_fin_req,
      return_mack => releaseLock_fin_ack,
      call_mdata => releaseLock_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseLock_instance:releaseLock-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => releaseLock_tag,
      lock_address_pointer => releaseLock_lock_address_pointer,
      start_req => releaseLock_start_req,
      start_ack => releaseLock_start_ack,
      fin_req => releaseLock_fin_req,
      fin_ack => releaseLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryByte_call_reqs => accessMemoryByte_call_reqs(0 downto 0),
      accessMemoryByte_call_acks => accessMemoryByte_call_acks(0 downto 0),
      accessMemoryByte_call_data => accessMemoryByte_call_data(144 downto 0),
      accessMemoryByte_call_tag => accessMemoryByte_call_tag(0 downto 0),
      accessMemoryByte_return_reqs => accessMemoryByte_return_reqs(0 downto 0),
      accessMemoryByte_return_acks => accessMemoryByte_return_acks(0 downto 0),
      accessMemoryByte_return_data => accessMemoryByte_return_data(7 downto 0),
      accessMemoryByte_return_tag => accessMemoryByte_return_tag(0 downto 0),
      tag_in => releaseLock_tag_in,
      tag_out => releaseLock_tag_out-- 
    ); -- 
  -- module setGlobalSignals
  -- call arbiter for module setGlobalSignals
  setGlobalSignals_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setGlobalSignals_call_reqs,
      call_acks => setGlobalSignals_call_acks,
      return_reqs => setGlobalSignals_return_reqs,
      return_acks => setGlobalSignals_return_acks,
      call_tag  => setGlobalSignals_call_tag,
      return_tag  => setGlobalSignals_return_tag,
      call_mtag => setGlobalSignals_tag_in,
      return_mtag => setGlobalSignals_tag_out,
      call_mreq => setGlobalSignals_start_req,
      call_mack => setGlobalSignals_start_ack,
      return_mreq => setGlobalSignals_fin_req,
      return_mack => setGlobalSignals_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  setGlobalSignals_instance:setGlobalSignals-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => setGlobalSignals_start_req,
      start_ack => setGlobalSignals_start_ack,
      fin_req => setGlobalSignals_fin_req,
      fin_ack => setGlobalSignals_fin_ack,
      clk => clk,
      reset => reset,
      NIC_INTR_ENABLE => NIC_INTR_ENABLE,
      NIC_INTR_INTERNAL => NIC_INTR_INTERNAL,
      NIC_INTR_pipe_write_req => NIC_INTR_pipe_write_req(1 downto 1),
      NIC_INTR_pipe_write_ack => NIC_INTR_pipe_write_ack(1 downto 1),
      NIC_INTR_pipe_write_data => NIC_INTR_pipe_write_data(1 downto 1),
      NIC_INTR_ENABLE_pipe_write_req => NIC_INTR_ENABLE_pipe_write_req(1 downto 1),
      NIC_INTR_ENABLE_pipe_write_ack => NIC_INTR_ENABLE_pipe_write_ack(1 downto 1),
      NIC_INTR_ENABLE_pipe_write_data => NIC_INTR_ENABLE_pipe_write_data(1 downto 1),
      MAC_ENABLE_pipe_write_req => MAC_ENABLE_pipe_write_req(1 downto 1),
      MAC_ENABLE_pipe_write_ack => MAC_ENABLE_pipe_write_ack(1 downto 1),
      MAC_ENABLE_pipe_write_data => MAC_ENABLE_pipe_write_data(1 downto 1),
      S_CONTROL_REGISTER_pipe_write_req => S_CONTROL_REGISTER_pipe_write_req(1 downto 1),
      S_CONTROL_REGISTER_pipe_write_ack => S_CONTROL_REGISTER_pipe_write_ack(1 downto 1),
      S_CONTROL_REGISTER_pipe_write_data => S_CONTROL_REGISTER_pipe_write_data(63 downto 32),
      S_NUMBER_OF_SERVERS_pipe_write_req => S_NUMBER_OF_SERVERS_pipe_write_req(1 downto 1),
      S_NUMBER_OF_SERVERS_pipe_write_ack => S_NUMBER_OF_SERVERS_pipe_write_ack(1 downto 1),
      S_NUMBER_OF_SERVERS_pipe_write_data => S_NUMBER_OF_SERVERS_pipe_write_data(63 downto 32),
      accessRegister_call_reqs => accessRegister_call_reqs(4 downto 4),
      accessRegister_call_acks => accessRegister_call_acks(4 downto 4),
      accessRegister_call_data => accessRegister_call_data(224 downto 180),
      accessRegister_call_tag => accessRegister_call_tag(9 downto 8),
      accessRegister_return_reqs => accessRegister_return_reqs(4 downto 4),
      accessRegister_return_acks => accessRegister_return_acks(4 downto 4),
      accessRegister_return_data => accessRegister_return_data(159 downto 128),
      accessRegister_return_tag => accessRegister_return_tag(9 downto 8),
      tag_in => setGlobalSignals_tag_in,
      tag_out => setGlobalSignals_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_tag <= setQueueElement_in_args(167 downto 160);
  setQueueElement_buf_base_address <= setQueueElement_in_args(159 downto 96);
  setQueueElement_write_index <= setQueueElement_in_args(95 downto 64);
  setQueueElement_q_w_data <= setQueueElement_in_args(63 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 168,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => setQueueElement_tag,
      buf_base_address => setQueueElement_buf_base_address,
      write_index => setQueueElement_write_index,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueElement_call_reqs => accessQueueElement_call_reqs(0 downto 0),
      accessQueueElement_call_acks => accessQueueElement_call_acks(0 downto 0),
      accessQueueElement_call_data => accessQueueElement_call_data(168 downto 0),
      accessQueueElement_call_tag => accessQueueElement_call_tag(0 downto 0),
      accessQueueElement_return_reqs => accessQueueElement_return_reqs(0 downto 0),
      accessQueueElement_return_acks => accessQueueElement_return_acks(0 downto 0),
      accessQueueElement_return_data => accessQueueElement_return_data(63 downto 0),
      accessQueueElement_return_tag => accessQueueElement_return_tag(0 downto 0),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_tag <= setQueuePointers_in_args(135 downto 128);
  setQueuePointers_q_base_address <= setQueuePointers_in_args(127 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 136,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => setQueuePointers_tag,
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueReadIndex_call_reqs => accessQueueReadIndex_call_reqs(1 downto 1),
      accessQueueReadIndex_call_acks => accessQueueReadIndex_call_acks(1 downto 1),
      accessQueueReadIndex_call_data => accessQueueReadIndex_call_data(209 downto 105),
      accessQueueReadIndex_call_tag => accessQueueReadIndex_call_tag(1 downto 1),
      accessQueueReadIndex_return_reqs => accessQueueReadIndex_return_reqs(1 downto 1),
      accessQueueReadIndex_return_acks => accessQueueReadIndex_return_acks(1 downto 1),
      accessQueueReadIndex_return_data => accessQueueReadIndex_return_data(63 downto 32),
      accessQueueReadIndex_return_tag => accessQueueReadIndex_return_tag(1 downto 1),
      accessQueueWriteIndex_call_reqs => accessQueueWriteIndex_call_reqs(1 downto 1),
      accessQueueWriteIndex_call_acks => accessQueueWriteIndex_call_acks(1 downto 1),
      accessQueueWriteIndex_call_data => accessQueueWriteIndex_call_data(209 downto 105),
      accessQueueWriteIndex_call_tag => accessQueueWriteIndex_call_tag(1 downto 1),
      accessQueueWriteIndex_return_reqs => accessQueueWriteIndex_return_reqs(1 downto 1),
      accessQueueWriteIndex_return_acks => accessQueueWriteIndex_return_acks(1 downto 1),
      accessQueueWriteIndex_return_data => accessQueueWriteIndex_return_data(63 downto 32),
      accessQueueWriteIndex_return_tag => accessQueueWriteIndex_return_tag(1 downto 1),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module setTotalMessages
  setTotalMessages_tag <= setTotalMessages_in_args(103 downto 96);
  setTotalMessages_q_base_address <= setTotalMessages_in_args(95 downto 32);
  setTotalMessages_updated_total_msgs <= setTotalMessages_in_args(31 downto 0);
  -- call arbiter for module setTotalMessages
  setTotalMessages_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 104,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setTotalMessages_call_reqs,
      call_acks => setTotalMessages_call_acks,
      return_reqs => setTotalMessages_return_reqs,
      return_acks => setTotalMessages_return_acks,
      call_data  => setTotalMessages_call_data,
      call_tag  => setTotalMessages_call_tag,
      return_tag  => setTotalMessages_return_tag,
      call_mtag => setTotalMessages_tag_in,
      return_mtag => setTotalMessages_tag_out,
      call_mreq => setTotalMessages_start_req,
      call_mack => setTotalMessages_start_ack,
      return_mreq => setTotalMessages_fin_req,
      return_mack => setTotalMessages_fin_ack,
      call_mdata => setTotalMessages_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setTotalMessages_instance:setTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      tag => setTotalMessages_tag,
      q_base_address => setTotalMessages_q_base_address,
      updated_total_msgs => setTotalMessages_updated_total_msgs,
      start_req => setTotalMessages_start_req,
      start_ack => setTotalMessages_start_ack,
      fin_req => setTotalMessages_fin_req,
      fin_ack => setTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessQueueTotalMsgs_call_reqs => accessQueueTotalMsgs_call_reqs(1 downto 1),
      accessQueueTotalMsgs_call_acks => accessQueueTotalMsgs_call_acks(1 downto 1),
      accessQueueTotalMsgs_call_data => accessQueueTotalMsgs_call_data(209 downto 105),
      accessQueueTotalMsgs_call_tag => accessQueueTotalMsgs_call_tag(1 downto 1),
      accessQueueTotalMsgs_return_reqs => accessQueueTotalMsgs_return_reqs(1 downto 1),
      accessQueueTotalMsgs_return_acks => accessQueueTotalMsgs_return_acks(1 downto 1),
      accessQueueTotalMsgs_return_data => accessQueueTotalMsgs_return_data(63 downto 32),
      accessQueueTotalMsgs_return_tag => accessQueueTotalMsgs_return_tag(1 downto 1),
      tag_in => setTotalMessages_tag_in,
      tag_out => setTotalMessages_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      S_CONTROL_REGISTER => S_CONTROL_REGISTER,
      S_NUMBER_OF_SERVERS => S_NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(15 downto 0),
      TX_ACTIVITY_LOGGER_pipe_write_req => TX_ACTIVITY_LOGGER_pipe_write_req(0 downto 0),
      TX_ACTIVITY_LOGGER_pipe_write_ack => TX_ACTIVITY_LOGGER_pipe_write_ack(0 downto 0),
      TX_ACTIVITY_LOGGER_pipe_write_data => TX_ACTIVITY_LOGGER_pipe_write_data(7 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(81 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(15 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(64 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      incrementNumberOfPacketsTransmitted_call_reqs => incrementNumberOfPacketsTransmitted_call_reqs(0 downto 0),
      incrementNumberOfPacketsTransmitted_call_acks => incrementNumberOfPacketsTransmitted_call_acks(0 downto 0),
      incrementNumberOfPacketsTransmitted_call_tag => incrementNumberOfPacketsTransmitted_call_tag(0 downto 0),
      incrementNumberOfPacketsTransmitted_return_reqs => incrementNumberOfPacketsTransmitted_return_reqs(0 downto 0),
      incrementNumberOfPacketsTransmitted_return_acks => incrementNumberOfPacketsTransmitted_return_acks(0 downto 0),
      incrementNumberOfPacketsTransmitted_return_tag => incrementNumberOfPacketsTransmitted_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(71 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_tag <= transmitPacket_in_args(71 downto 64);
  transmitPacket_packet_pointer <= transmitPacket_in_args(63 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => transmitPacket_tag,
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 0),
      accessMemoryDword_call_reqs => accessMemoryDword_call_reqs(1 downto 0),
      accessMemoryDword_call_acks => accessMemoryDword_call_acks(1 downto 0),
      accessMemoryDword_call_data => accessMemoryDword_call_data(401 downto 0),
      accessMemoryDword_call_tag => accessMemoryDword_call_tag(3 downto 0),
      accessMemoryDword_return_reqs => accessMemoryDword_return_reqs(1 downto 0),
      accessMemoryDword_return_acks => accessMemoryDword_return_acks(1 downto 0),
      accessMemoryDword_return_data => accessMemoryDword_return_data(127 downto 0),
      accessMemoryDword_return_tag => accessMemoryDword_return_tag(3 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_tag <= writeControlInformationToMem_in_args(106 downto 99);
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(98 downto 35);
  writeControlInformationToMem_max_addr_offset <= writeControlInformationToMem_in_args(34 downto 19);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(18 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 107,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => writeControlInformationToMem_tag,
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      max_addr_offset => writeControlInformationToMem_max_addr_offset,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemoryDword_call_reqs => accessMemoryDword_call_reqs(3 downto 3),
      accessMemoryDword_call_acks => accessMemoryDword_call_acks(3 downto 3),
      accessMemoryDword_call_data => accessMemoryDword_call_data(803 downto 603),
      accessMemoryDword_call_tag => accessMemoryDword_call_tag(7 downto 6),
      accessMemoryDword_return_reqs => accessMemoryDword_return_reqs(3 downto 3),
      accessMemoryDword_return_acks => accessMemoryDword_return_acks(3 downto 3),
      accessMemoryDword_return_data => accessMemoryDword_return_data(255 downto 192),
      accessMemoryDword_return_tag => accessMemoryDword_return_tag(7 downto 6),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_tag <= writeEthernetHeaderToMem_in_args(71 downto 64);
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(63 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_addr_offset ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => writeEthernetHeaderToMem_tag,
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      addr_offset => writeEthernetHeaderToMem_addr_offset,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemoryDword_call_reqs => accessMemoryDword_call_reqs(6 downto 6),
      accessMemoryDword_call_acks => accessMemoryDword_call_acks(6 downto 6),
      accessMemoryDword_call_data => accessMemoryDword_call_data(1406 downto 1206),
      accessMemoryDword_call_tag => accessMemoryDword_call_tag(13 downto 12),
      accessMemoryDword_return_reqs => accessMemoryDword_return_reqs(6 downto 6),
      accessMemoryDword_return_acks => accessMemoryDword_return_acks(6 downto 6),
      accessMemoryDword_return_data => accessMemoryDword_return_data(447 downto 384),
      accessMemoryDword_return_tag => accessMemoryDword_return_tag(13 downto 12),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_tag <= writePayloadToMem_in_args(103 downto 96);
  writePayloadToMem_max_addr_offset <= writePayloadToMem_in_args(95 downto 80);
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(79 downto 16);
  writePayloadToMem_addr_offset <= writePayloadToMem_in_args(15 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_11 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 104,
      return_data_width => 20,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      tag => writePayloadToMem_tag,
      max_addr_offset => writePayloadToMem_max_addr_offset,
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      addr_offset => writePayloadToMem_addr_offset,
      packet_size_11 => writePayloadToMem_packet_size_11,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemoryDword_call_reqs => accessMemoryDword_call_reqs(4 downto 4),
      accessMemoryDword_call_acks => accessMemoryDword_call_acks(4 downto 4),
      accessMemoryDword_call_data => accessMemoryDword_call_data(1004 downto 804),
      accessMemoryDword_call_tag => accessMemoryDword_call_tag(9 downto 8),
      accessMemoryDword_return_reqs => accessMemoryDword_return_reqs(4 downto 4),
      accessMemoryDword_return_acks => accessMemoryDword_return_acks(4 downto 4),
      accessMemoryDword_return_data => accessMemoryDword_return_data(319 downto 256),
      accessMemoryDword_return_tag => accessMemoryDword_return_tag(9 downto 8),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 8 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 8 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MAC_ENABLE_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe MAC_ENABLE",
      volatile_flag => false,
      num_writes => 2,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => MAC_ENABLE,
      write_req => MAC_ENABLE_pipe_write_req,
      write_ack => MAC_ENABLE_pipe_write_ack,
      write_data => MAC_ENABLE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_DEBUG_SIGNAL_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NIC_DEBUG_SIGNAL",
      volatile_flag => false,
      num_writes => 1,
      data_width => 256 --
    ) 
    port map( -- 
      read_data => NIC_DEBUG_SIGNAL,
      write_req => NIC_DEBUG_SIGNAL_pipe_write_req,
      write_ack => NIC_DEBUG_SIGNAL_pipe_write_ack,
      write_data => NIC_DEBUG_SIGNAL_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_INTR_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NIC_INTR",
      volatile_flag => false,
      num_writes => 2,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => NIC_INTR,
      write_req => NIC_INTR_pipe_write_req,
      write_ack => NIC_INTR_pipe_write_ack,
      write_data => NIC_INTR_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_INTR_ENABLE_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NIC_INTR_ENABLE",
      volatile_flag => false,
      num_writes => 2,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => NIC_INTR_ENABLE,
      write_req => NIC_INTR_ENABLE_pipe_write_req,
      write_ack => NIC_INTR_ENABLE_pipe_write_ack,
      write_data => NIC_INTR_ENABLE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_INTR_INTERNAL_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NIC_INTR_INTERNAL",
      volatile_flag => false,
      num_writes => 1,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => NIC_INTR_INTERNAL,
      write_req => NIC_INTR_INTERNAL_pipe_write_req,
      write_ack => NIC_INTR_INTERNAL_pipe_write_ack,
      write_data => NIC_INTR_INTERNAL_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  QUEUE_MONITOR_SIGNAL_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe QUEUE_MONITOR_SIGNAL",
      volatile_flag => false,
      num_writes => 2,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => QUEUE_MONITOR_SIGNAL,
      write_req => QUEUE_MONITOR_SIGNAL_pipe_write_req,
      write_ack => QUEUE_MONITOR_SIGNAL_pipe_write_ack,
      write_data => QUEUE_MONITOR_SIGNAL_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  RX_ACTIVITY_LOGGER_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe RX_ACTIVITY_LOGGER",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => RX_ACTIVITY_LOGGER_pipe_read_req,
      read_ack => RX_ACTIVITY_LOGGER_pipe_read_ack,
      read_data => RX_ACTIVITY_LOGGER_pipe_read_data,
      write_req => RX_ACTIVITY_LOGGER_pipe_write_req,
      write_ack => RX_ACTIVITY_LOGGER_pipe_write_ack,
      write_data => RX_ACTIVITY_LOGGER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  S_CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe S_CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 2,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => S_CONTROL_REGISTER,
      write_req => S_CONTROL_REGISTER_pipe_write_req,
      write_ack => S_CONTROL_REGISTER_pipe_write_ack,
      write_data => S_CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  S_NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe S_NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 2,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => S_NUMBER_OF_SERVERS,
      write_req => S_NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => S_NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => S_NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  TX_ACTIVITY_LOGGER_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe TX_ACTIVITY_LOGGER",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => TX_ACTIVITY_LOGGER_pipe_read_req,
      read_ack => TX_ACTIVITY_LOGGER_pipe_read_ack,
      read_data => TX_ACTIVITY_LOGGER_pipe_read_data,
      write_req => TX_ACTIVITY_LOGGER_pipe_write_req,
      write_ack => TX_ACTIVITY_LOGGER_pipe_write_ack,
      write_data => TX_ACTIVITY_LOGGER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  memory_access_lock_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe memory_access_lock",
      num_reads => 1,
      num_writes => 2,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => memory_access_lock_pipe_read_req,
      read_ack => memory_access_lock_pipe_read_ack,
      read_data => memory_access_lock_pipe_read_data,
      write_req => memory_access_lock_pipe_write_req,
      write_ack => memory_access_lock_pipe_write_ack,
      write_data => memory_access_lock_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end nic_arch;

-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity AccessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    register_index : in  std_logic_vector(5 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity AccessRegister;
architecture AccessRegister_arch of AccessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal register_index_buffer :  std_logic_vector(5 downto 0);
  signal register_index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal AccessRegister_CP_0_start: Boolean;
  signal AccessRegister_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_req_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_req_1 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_ack_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_req_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_ack_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_req_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "AccessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(10 downto 5) <= register_index;
  register_index_buffer <= in_buffer_data_out(10 downto 5);
  in_buffer_data_in(42 downto 11) <= wdata;
  wdata_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  AccessRegister_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "AccessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  AccessRegister_CP_0: Block -- control-path 
    signal AccessRegister_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    AccessRegister_CP_0_elements(0) <= AccessRegister_CP_0_start;
    AccessRegister_CP_0_symbol <= AccessRegister_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_sample_start_
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Sample/req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/$entry
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_sample_start_
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_sample_completed_
      -- CP-element group 1: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_update_start_
      -- CP-element group 1: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Sample/ack
      -- CP-element group 1: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Update/$entry
      -- CP-element group 1: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_ack_0, ack => AccessRegister_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(1), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_update_completed_
      -- CP-element group 2: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Update/$exit
      -- CP-element group 2: 	 assign_stmt_82_to_assign_stmt_100/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_ack_1, ack => AccessRegister_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_sample_completed_
      -- CP-element group 3: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_update_start_
      -- CP-element group 3: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Sample/ra
      -- CP-element group 3: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Update/$entry
      -- CP-element group 3: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_ack_0, ack => AccessRegister_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(3), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_update_completed_
      -- CP-element group 4: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Update/$exit
      -- CP-element group 4: 	 assign_stmt_82_to_assign_stmt_100/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_ack_1, ack => AccessRegister_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_82_to_assign_stmt_100/$exit
      -- 
    AccessRegister_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "AccessRegister_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= AccessRegister_CP_0_elements(4) & AccessRegister_CP_0_elements(2);
      gj_AccessRegister_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => AccessRegister_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_77_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u6_u38_80_wire : std_logic_vector(37 downto 0);
    signal request_82 : std_logic_vector(42 downto 0);
    signal response_94 : std_logic_vector(32 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_99_inst
    rdata_buffer <= response_94(31 downto 0);
    -- binary operator CONCAT_u1_u5_77_inst
    process(rwbar_buffer, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(rwbar_buffer, bmask_buffer, tmp_var);
      CONCAT_u1_u5_77_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u5_u43_81_inst
    process(CONCAT_u1_u5_77_wire, CONCAT_u6_u38_80_wire) -- 
      variable tmp_var : std_logic_vector(42 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_77_wire, CONCAT_u6_u38_80_wire, tmp_var);
      request_82 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u38_80_inst
    process(register_index_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(register_index_buffer, wdata_buffer, tmp_var);
      CONCAT_u6_u38_80_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_req_0;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_req_1;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_93_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_94 <= data_out(32 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_req_0;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_req_1;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_88_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_82;
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE", data_width => 43, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end AccessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity NicRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
    MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity NicRegisterAccessDaemon;
architecture NicRegisterAccessDaemon_arch of NicRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal NicRegisterAccessDaemon_CP_116_start: Boolean;
  signal NicRegisterAccessDaemon_CP_116_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal array_obj_ref_193_store_0_req_0 : boolean;
  signal array_obj_ref_193_store_0_ack_0 : boolean;
  signal array_obj_ref_193_store_0_req_1 : boolean;
  signal array_obj_ref_193_store_0_ack_1 : boolean;
  signal MUX_208_inst_req_0 : boolean;
  signal MUX_208_inst_ack_0 : boolean;
  signal MUX_208_inst_req_1 : boolean;
  signal MUX_208_inst_ack_1 : boolean;
  signal WPIPE_MAC_ENABLE_202_inst_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_202_inst_ack_0 : boolean;
  signal WPIPE_MAC_ENABLE_202_inst_req_1 : boolean;
  signal WPIPE_MAC_ENABLE_202_inst_ack_1 : boolean;
  signal if_stmt_210_branch_req_0 : boolean;
  signal if_stmt_210_branch_ack_1 : boolean;
  signal if_stmt_210_branch_ack_0 : boolean;
  signal phi_stmt_185_req_0 : boolean;
  signal nI_201_190_buf_req_0 : boolean;
  signal nI_201_190_buf_ack_0 : boolean;
  signal nI_201_190_buf_req_1 : boolean;
  signal nI_201_190_buf_ack_1 : boolean;
  signal phi_stmt_185_req_1 : boolean;
  signal phi_stmt_185_ack_0 : boolean;
  signal do_while_stmt_219_branch_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_ack_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_req_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_ack_1 : boolean;
  signal array_obj_ref_243_load_0_req_0 : boolean;
  signal array_obj_ref_243_load_0_ack_0 : boolean;
  signal array_obj_ref_243_load_0_req_1 : boolean;
  signal array_obj_ref_243_load_0_ack_1 : boolean;
  signal W_rwbar_252_delayed_5_0_248_inst_req_0 : boolean;
  signal W_rwbar_252_delayed_5_0_248_inst_ack_0 : boolean;
  signal W_rwbar_252_delayed_5_0_248_inst_req_1 : boolean;
  signal W_rwbar_252_delayed_5_0_248_inst_ack_1 : boolean;
  signal W_bmask_253_delayed_5_0_251_inst_req_0 : boolean;
  signal W_bmask_253_delayed_5_0_251_inst_ack_0 : boolean;
  signal W_bmask_253_delayed_5_0_251_inst_req_1 : boolean;
  signal W_bmask_253_delayed_5_0_251_inst_ack_1 : boolean;
  signal W_wdata_255_delayed_5_0_254_inst_req_0 : boolean;
  signal W_wdata_255_delayed_5_0_254_inst_ack_0 : boolean;
  signal W_wdata_255_delayed_5_0_254_inst_req_1 : boolean;
  signal W_wdata_255_delayed_5_0_254_inst_ack_1 : boolean;
  signal W_index_256_delayed_5_0_257_inst_req_0 : boolean;
  signal W_index_256_delayed_5_0_257_inst_ack_0 : boolean;
  signal W_index_256_delayed_5_0_257_inst_req_1 : boolean;
  signal W_index_256_delayed_5_0_257_inst_ack_1 : boolean;
  signal call_stmt_266_call_req_0 : boolean;
  signal call_stmt_266_call_ack_0 : boolean;
  signal call_stmt_266_call_req_1 : boolean;
  signal call_stmt_266_call_ack_1 : boolean;
  signal W_rwbar_260_delayed_5_0_267_inst_req_0 : boolean;
  signal W_rwbar_260_delayed_5_0_267_inst_ack_0 : boolean;
  signal W_rwbar_260_delayed_5_0_267_inst_req_1 : boolean;
  signal W_rwbar_260_delayed_5_0_267_inst_ack_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_req_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_ack_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_req_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_ack_1 : boolean;
  signal do_while_stmt_219_branch_ack_0 : boolean;
  signal do_while_stmt_219_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  NicRegisterAccessDaemon_CP_116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  NicRegisterAccessDaemon_CP_116: Block -- control-path 
    signal NicRegisterAccessDaemon_CP_116_elements: BooleanArray(65 downto 0);
    -- 
  begin -- 
    NicRegisterAccessDaemon_CP_116_elements(0) <= NicRegisterAccessDaemon_CP_116_start;
    NicRegisterAccessDaemon_CP_116_symbol <= NicRegisterAccessDaemon_CP_116_elements(16);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_183/$entry
      -- CP-element group 0: 	 branch_block_stmt_183/branch_block_stmt_183__entry__
      -- CP-element group 0: 	 branch_block_stmt_183/merge_stmt_184__entry__
      -- CP-element group 0: 	 branch_block_stmt_183/merge_stmt_184_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/phi_stmt_185/$entry
      -- CP-element group 0: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/phi_stmt_185/phi_stmt_185_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	15 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_sample_completed_
      -- 
    ra_183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_193_store_0_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	15 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/word_access_complete/word_0/ca
      -- 
    ca_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_193_store_0_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_start/ack
      -- 
    ack_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_208_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_complete/ack
      -- CP-element group 4: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Sample/req
      -- 
    ack_208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_208_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(4)); -- 
    req_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(4), ack => WPIPE_MAC_ENABLE_202_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_update_start_
      -- CP-element group 5: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Update/req
      -- 
    ack_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_202_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(5)); -- 
    req_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(5), ack => WPIPE_MAC_ENABLE_202_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/WPIPE_MAC_ENABLE_202_Update/ack
      -- 
    ack_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_202_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(6)); -- 
    -- CP-element group 7:  branch  join  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (24) 
      -- CP-element group 7: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209__exit__
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210__entry__
      -- CP-element group 7: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_dead_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/ULT_u7_u1_213_inputs/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/ULT_u7_u1_213_inputs/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/ULT_u7_u1_213/SplitProtocol/Update/ca
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_eval_test/branch_req
      -- CP-element group 7: 	 branch_block_stmt_183/ULT_u7_u1_213_place
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_if_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_183/if_stmt_210_else_link/$entry
      -- 
    branch_req_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(7), ack => if_stmt_210_branch_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 42) := "NicRegisterAccessDaemon_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(2) & NicRegisterAccessDaemon_CP_116_elements(6);
      gj_NicRegisterAccessDaemon_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	12 
    -- CP-element group 8:  members (11) 
      -- CP-element group 8: 	 branch_block_stmt_183/if_stmt_210_if_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_183/if_stmt_210_if_link/if_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_183/loopback
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/$entry
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/$entry
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Sample/req
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Update/req
      -- 
    if_choice_transition_254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_210_branch_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(8)); -- 
    req_290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(8), ack => nI_201_190_buf_req_0); -- 
    req_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(8), ack => nI_201_190_buf_req_1); -- 
    -- CP-element group 9:  merge  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	17 
    -- CP-element group 9:  members (8) 
      -- CP-element group 9: 	 branch_block_stmt_183/$exit
      -- CP-element group 9: 	 branch_block_stmt_183/branch_block_stmt_183__exit__
      -- CP-element group 9: 	 branch_block_stmt_183/if_stmt_210__exit__
      -- CP-element group 9: 	 branch_block_stmt_183/if_stmt_210_else_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_183/if_stmt_210_else_link/else_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_218/$entry
      -- CP-element group 9: 	 branch_block_stmt_218/branch_block_stmt_218__entry__
      -- CP-element group 9: 	 branch_block_stmt_218/do_while_stmt_219__entry__
      -- 
    else_choice_transition_258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_210_branch_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(9)); -- 
    -- CP-element group 10:  transition  output  delay-element  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	14 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/$exit
      -- CP-element group 10: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/phi_stmt_185/$exit
      -- CP-element group 10: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/phi_stmt_185/phi_stmt_185_sources/$exit
      -- CP-element group 10: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/phi_stmt_185/phi_stmt_185_sources/type_cast_189_konst_delay_trans
      -- CP-element group 10: 	 branch_block_stmt_183/merge_stmt_184__entry___PhiReq/phi_stmt_185/phi_stmt_185_req
      -- 
    phi_stmt_185_req_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_185_req_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(10), ack => phi_stmt_185_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(10) is a control-delay.
    cp_element_10_delay: control_delay_element  generic map(name => " 10_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(0), ack => NicRegisterAccessDaemon_CP_116_elements(10), clk => clk, reset =>reset);
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Sample/ack
      -- 
    ack_291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_201_190_buf_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/Update/ack
      -- 
    ack_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_201_190_buf_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_183/loopback_PhiReq/$exit
      -- CP-element group 13: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/$exit
      -- CP-element group 13: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/$exit
      -- CP-element group 13: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_sources/Interlock/$exit
      -- CP-element group 13: 	 branch_block_stmt_183/loopback_PhiReq/phi_stmt_185/phi_stmt_185_req
      -- 
    phi_stmt_185_req_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_185_req_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(13), ack => phi_stmt_185_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(11) & NicRegisterAccessDaemon_CP_116_elements(12);
      gj_NicRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  merge  transition  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: 	10 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_183/merge_stmt_184_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_183/merge_stmt_184_PhiAck/$entry
      -- 
    NicRegisterAccessDaemon_CP_116_elements(14) <= OrReduce(NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(10));
    -- CP-element group 15:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: 	1 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	3 
    -- CP-element group 15:  members (51) 
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/array_obj_ref_193_Split/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/array_obj_ref_193_Split/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/array_obj_ref_193_Split/split_req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/array_obj_ref_193_Split/split_ack
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_183/merge_stmt_184__exit__
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209__entry__
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_update_start_
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_final_index_sum_regn/req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/array_obj_ref_193_Update/word_access_complete/word_0/cr
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_update_start_
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_start/req
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_183/assign_stmt_196_to_assign_stmt_209/MUX_208_complete/req
      -- CP-element group 15: 	 branch_block_stmt_183/merge_stmt_184_PhiAck/$exit
      -- CP-element group 15: 	 branch_block_stmt_183/merge_stmt_184_PhiAck/phi_stmt_185_ack
      -- 
    phi_stmt_185_ack_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_185_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(15)); -- 
    rr_182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => array_obj_ref_193_store_0_req_0); -- 
    cr_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => array_obj_ref_193_store_0_req_1); -- 
    req_202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => MUX_208_inst_req_0); -- 
    req_207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => MUX_208_inst_req_1); -- 
    -- CP-element group 16:  transition  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	65 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (4) 
      -- CP-element group 16: 	 $exit
      -- CP-element group 16: 	 branch_block_stmt_218/$exit
      -- CP-element group 16: 	 branch_block_stmt_218/branch_block_stmt_218__exit__
      -- CP-element group 16: 	 branch_block_stmt_218/do_while_stmt_219__exit__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(16) <= NicRegisterAccessDaemon_CP_116_elements(65);
    -- CP-element group 17:  transition  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	23 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_218/do_while_stmt_219/$entry
      -- CP-element group 17: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219__entry__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(17) <= NicRegisterAccessDaemon_CP_116_elements(9);
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219__exit__
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(18) is bound as output of CP function.
    -- CP-element group 19:  merge  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_218/do_while_stmt_219/loop_back
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(19) is bound as output of CP function.
    -- CP-element group 20:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	60 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20: 	64 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_218/do_while_stmt_219/condition_done
      -- CP-element group 20: 	 branch_block_stmt_218/do_while_stmt_219/loop_exit/$entry
      -- CP-element group 20: 	 branch_block_stmt_218/do_while_stmt_219/loop_taken/$entry
      -- 
    NicRegisterAccessDaemon_CP_116_elements(20) <= NicRegisterAccessDaemon_CP_116_elements(60);
    -- CP-element group 21:  branch  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	62 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_218/do_while_stmt_219/loop_body_done
      -- 
    NicRegisterAccessDaemon_CP_116_elements(21) <= NicRegisterAccessDaemon_CP_116_elements(62);
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/back_edge_to_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(22) <= NicRegisterAccessDaemon_CP_116_elements(19);
    -- CP-element group 23:  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/first_time_through_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(23) <= NicRegisterAccessDaemon_CP_116_elements(17);
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	60 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/$entry
      -- CP-element group 24: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/loop_body_start
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Sample/rr
      -- 
    rr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(25), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(24) & NicRegisterAccessDaemon_CP_116_elements(28);
      gj_NicRegisterAccessDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	35 
    -- CP-element group 26: 	39 
    -- CP-element group 26: 	43 
    -- CP-element group 26: 	47 
    -- CP-element group 26: 	55 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_update_start_
      -- CP-element group 26: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Update/cr
      -- 
    cr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(26), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(27) & NicRegisterAccessDaemon_CP_116_elements(31) & NicRegisterAccessDaemon_CP_116_elements(35) & NicRegisterAccessDaemon_CP_116_elements(39) & NicRegisterAccessDaemon_CP_116_elements(43) & NicRegisterAccessDaemon_CP_116_elements(47) & NicRegisterAccessDaemon_CP_116_elements(55);
      gj_NicRegisterAccessDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Sample/ra
      -- 
    ra_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	33 
    -- CP-element group 28: 	37 
    -- CP-element group 28: 	41 
    -- CP-element group 28: 	45 
    -- CP-element group 28: 	53 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (29) 
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_word_address_calculated
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_root_address_calculated
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_offset_calculated
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_resized_0
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_scaled_0
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_computed_0
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_resize_0/$entry
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_resize_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_resize_0/index_resize_req
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_resize_0/index_resize_ack
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_scale_0/$entry
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_scale_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_scale_0/scale_rename_req
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_index_scale_0/scale_rename_ack
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_final_index_sum_regn/$entry
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_final_index_sum_regn/$exit
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_final_index_sum_regn/req
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_final_index_sum_regn/ack
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_base_plus_offset/$entry
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_base_plus_offset/$exit
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_word_addrgen/$entry
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_word_addrgen/$exit
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_word_addrgen/root_register_req
      -- CP-element group 28: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_word_addrgen/root_register_ack
      -- 
    ca_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: 	52 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/word_access_start/word_0/rr
      -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(29), ack => array_obj_ref_243_load_0_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(31) & NicRegisterAccessDaemon_CP_116_elements(52);
      gj_NicRegisterAccessDaemon_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	51 
    -- CP-element group 30: 	58 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_update_start_
      -- CP-element group 30: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/word_access_complete/$entry
      -- CP-element group 30: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/word_access_complete/word_0/$entry
      -- CP-element group 30: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/word_access_complete/word_0/cr
      -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(30), ack => array_obj_ref_243_load_0_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(32) & NicRegisterAccessDaemon_CP_116_elements(51) & NicRegisterAccessDaemon_CP_116_elements(58);
      gj_NicRegisterAccessDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	61 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Sample/word_access_start/word_0/ra
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_243_load_0_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	49 
    -- CP-element group 32: 	57 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/array_obj_ref_243_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/array_obj_ref_243_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/array_obj_ref_243_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_Update/array_obj_ref_243_Merge/merge_ack
      -- 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_243_load_0_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	28 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Sample/req
      -- 
    req_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(33), ack => W_rwbar_252_delayed_5_0_248_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(35);
      gj_NicRegisterAccessDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	51 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_update_start_
      -- CP-element group 34: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Update/req
      -- 
    req_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(34), ack => W_rwbar_252_delayed_5_0_248_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(36) & NicRegisterAccessDaemon_CP_116_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	26 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Sample/ack
      -- 
    ack_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_252_delayed_5_0_248_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	49 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_250_Update/ack
      -- 
    ack_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_252_delayed_5_0_248_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	28 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Sample/req
      -- 
    req_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(37), ack => W_bmask_253_delayed_5_0_251_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(39);
      gj_NicRegisterAccessDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: 	51 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_update_start_
      -- CP-element group 38: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Update/req
      -- 
    req_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(38), ack => W_bmask_253_delayed_5_0_251_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(40) & NicRegisterAccessDaemon_CP_116_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	26 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Sample/ack
      -- 
    ack_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_253_delayed_5_0_251_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_253_Update/ack
      -- 
    ack_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_253_delayed_5_0_251_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	28 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Sample/req
      -- 
    req_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(41), ack => W_wdata_255_delayed_5_0_254_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	51 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_update_start_
      -- CP-element group 42: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Update/req
      -- 
    req_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(42), ack => W_wdata_255_delayed_5_0_254_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(44) & NicRegisterAccessDaemon_CP_116_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	26 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Sample/ack
      -- 
    ack_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_255_delayed_5_0_254_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	49 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_256_Update/ack
      -- 
    ack_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_255_delayed_5_0_254_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	28 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Sample/req
      -- 
    req_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(45), ack => W_index_256_delayed_5_0_257_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(47);
      gj_NicRegisterAccessDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: 	51 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_update_start_
      -- CP-element group 46: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Update/req
      -- 
    req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(46), ack => W_index_256_delayed_5_0_257_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(48) & NicRegisterAccessDaemon_CP_116_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	26 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Sample/ack
      -- 
    ack_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_256_delayed_5_0_257_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(47)); -- 
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_259_Update/ack
      -- 
    ack_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_256_delayed_5_0_257_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	32 
    -- CP-element group 49: 	36 
    -- CP-element group 49: 	40 
    -- CP-element group 49: 	44 
    -- CP-element group 49: 	48 
    -- CP-element group 49: 	61 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Sample/crr
      -- 
    crr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(49), ack => call_stmt_266_call_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 31,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(32) & NicRegisterAccessDaemon_CP_116_elements(36) & NicRegisterAccessDaemon_CP_116_elements(40) & NicRegisterAccessDaemon_CP_116_elements(44) & NicRegisterAccessDaemon_CP_116_elements(48) & NicRegisterAccessDaemon_CP_116_elements(61) & NicRegisterAccessDaemon_CP_116_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_update_start_
      -- CP-element group 50: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Update/ccr
      -- 
    ccr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(50), ack => call_stmt_266_call_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(52);
      gj_NicRegisterAccessDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	30 
    -- CP-element group 51: 	34 
    -- CP-element group 51: 	38 
    -- CP-element group 51: 	42 
    -- CP-element group 51: 	46 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Sample/cra
      -- 
    cra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_266_call_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	62 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	29 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/call_stmt_266_Update/cca
      -- CP-element group 52: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/ring_reenable_memory_space_0
      -- 
    cca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_266_call_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	28 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Sample/req
      -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(53), ack => W_rwbar_260_delayed_5_0_267_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(55);
      gj_NicRegisterAccessDaemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	58 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_update_start_
      -- CP-element group 54: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Update/req
      -- 
    req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(54), ack => W_rwbar_260_delayed_5_0_267_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(56) & NicRegisterAccessDaemon_CP_116_elements(58);
      gj_NicRegisterAccessDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	26 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Sample/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_260_delayed_5_0_267_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/assign_stmt_269_Update/ack
      -- 
    ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_260_delayed_5_0_267_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	56 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Sample/req
      -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(57), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(32) & NicRegisterAccessDaemon_CP_116_elements(56) & NicRegisterAccessDaemon_CP_116_elements(59);
      gj_NicRegisterAccessDaemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	30 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_update_start_
      -- CP-element group 58: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Update/req
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(58)); -- 
    req_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(58), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	62 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_Update/ack
      -- 
    ack_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(59)); -- 
    -- CP-element group 60:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	24 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	20 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/condition_evaluated
      -- CP-element group 60: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(60), ack => do_while_stmt_219_branch_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(24), ack => NicRegisterAccessDaemon_CP_116_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	31 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	49 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/array_obj_ref_243_call_stmt_266_delay
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(61) is a control-delay.
    cp_element_61_delay: control_delay_element  generic map(name => " 61_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(31), ack => NicRegisterAccessDaemon_CP_116_elements(61), clk => clk, reset =>reset);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	52 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	21 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_218/do_while_stmt_219/do_while_stmt_219_loop_body/$exit
      -- 
    NicRegisterAccessDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(52) & NicRegisterAccessDaemon_CP_116_elements(59);
      gj_NicRegisterAccessDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_218/do_while_stmt_219/loop_exit/$exit
      -- CP-element group 63: 	 branch_block_stmt_218/do_while_stmt_219/loop_exit/ack
      -- 
    ack_507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_219_branch_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	20 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_218/do_while_stmt_219/loop_taken/$exit
      -- CP-element group 64: 	 branch_block_stmt_218/do_while_stmt_219/loop_taken/ack
      -- 
    ack_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_219_branch_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(64)); -- 
    -- CP-element group 65:  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	16 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_218/do_while_stmt_219/$exit
      -- 
    NicRegisterAccessDaemon_CP_116_elements(65) <= NicRegisterAccessDaemon_CP_116_elements(18);
    NicRegisterAccessDaemon_do_while_stmt_219_terminator_512: loop_terminator -- 
      generic map (name => " NicRegisterAccessDaemon_do_while_stmt_219_terminator_512", max_iterations_in_flight =>31) 
      port map(loop_body_exit => NicRegisterAccessDaemon_CP_116_elements(21),loop_continue => NicRegisterAccessDaemon_CP_116_elements(64),loop_terminate => NicRegisterAccessDaemon_CP_116_elements(63),loop_back => NicRegisterAccessDaemon_CP_116_elements(19),loop_exit => NicRegisterAccessDaemon_CP_116_elements(18),clk => clk, reset => reset); -- 
    entry_tmerge_325_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= NicRegisterAccessDaemon_CP_116_elements(22);
        preds(1)  <= NicRegisterAccessDaemon_CP_116_elements(23);
        entry_tmerge_325 : transition_merge -- 
          generic map(name => " entry_tmerge_325")
          port map (preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(24));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u7_u1_205_wire : std_logic_vector(0 downto 0);
    signal I_185 : std_logic_vector(6 downto 0);
    signal MUX_208_wire : std_logic_vector(0 downto 0);
    signal R_I_192_resized : std_logic_vector(5 downto 0);
    signal R_I_192_scaled : std_logic_vector(5 downto 0);
    signal R_index_242_resized : std_logic_vector(5 downto 0);
    signal R_index_242_scaled : std_logic_vector(5 downto 0);
    signal ULT_u7_u1_213_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_193_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_193_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_193_word_offset_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_243_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_243_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_243_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_243_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_243_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_243_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_243_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_232 : std_logic_vector(3 downto 0);
    signal bmask_253_delayed_5_0_253 : std_logic_vector(3 downto 0);
    signal index_236 : std_logic_vector(5 downto 0);
    signal index_256_delayed_5_0_259 : std_logic_vector(5 downto 0);
    signal konst_199_wire_constant : std_logic_vector(6 downto 0);
    signal konst_204_wire_constant : std_logic_vector(6 downto 0);
    signal konst_206_wire_constant : std_logic_vector(0 downto 0);
    signal konst_207_wire_constant : std_logic_vector(0 downto 0);
    signal konst_212_wire_constant : std_logic_vector(6 downto 0);
    signal konst_287_wire_constant : std_logic_vector(0 downto 0);
    signal nI_201 : std_logic_vector(6 downto 0);
    signal nI_201_190_buffered : std_logic_vector(6 downto 0);
    signal rdata_276 : std_logic_vector(31 downto 0);
    signal req_223 : std_logic_vector(42 downto 0);
    signal resp_282 : std_logic_vector(32 downto 0);
    signal rval_244 : std_logic_vector(31 downto 0);
    signal rwbar_228 : std_logic_vector(0 downto 0);
    signal rwbar_252_delayed_5_0_250 : std_logic_vector(0 downto 0);
    signal rwbar_260_delayed_5_0_269 : std_logic_vector(0 downto 0);
    signal type_cast_189_wire_constant : std_logic_vector(6 downto 0);
    signal type_cast_195_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_274_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_279_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_240 : std_logic_vector(31 downto 0);
    signal wdata_255_delayed_5_0_256 : std_logic_vector(31 downto 0);
    signal wval_266 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_193_offset_scale_factor_0 <= "000001";
    array_obj_ref_193_resized_base_address <= "000000";
    array_obj_ref_193_word_offset_0 <= "000000";
    array_obj_ref_243_offset_scale_factor_0 <= "000001";
    array_obj_ref_243_resized_base_address <= "000000";
    array_obj_ref_243_word_offset_0 <= "000000";
    konst_199_wire_constant <= "0000001";
    konst_204_wire_constant <= "0111111";
    konst_206_wire_constant <= "1";
    konst_207_wire_constant <= "0";
    konst_212_wire_constant <= "0111111";
    konst_287_wire_constant <= "1";
    type_cast_189_wire_constant <= "0000000";
    type_cast_195_wire_constant <= "00000000000000000000000000000000";
    type_cast_274_wire_constant <= "00000000000000000000000000000000";
    type_cast_279_wire_constant <= "0";
    phi_stmt_185: Block -- phi operator 
      signal idata: std_logic_vector(13 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_189_wire_constant & nI_201_190_buffered;
      req <= phi_stmt_185_req_0 & phi_stmt_185_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_185",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 7) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_185_ack_0,
          idata => idata,
          odata => I_185,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_185
    MUX_208_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_208_inst_req_0;
      MUX_208_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_208_inst_req_1;
      MUX_208_inst_ack_1<= update_ack(0);
      MUX_208_inst: SelectSplitProtocol generic map(name => "MUX_208_inst", data_width => 1, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => konst_206_wire_constant, y => konst_207_wire_constant, sel => EQ_u7_u1_205_wire, z => MUX_208_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_275_inst
    rdata_276 <= rval_244 when (rwbar_260_delayed_5_0_269(0) /=  '0') else type_cast_274_wire_constant;
    -- flow-through slice operator slice_227_inst
    rwbar_228 <= req_223(42 downto 42);
    -- flow-through slice operator slice_231_inst
    bmask_232 <= req_223(41 downto 38);
    -- flow-through slice operator slice_235_inst
    index_236 <= req_223(37 downto 32);
    -- flow-through slice operator slice_239_inst
    wdata_240 <= req_223(31 downto 0);
    W_bmask_253_delayed_5_0_251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_253_delayed_5_0_251_inst_req_0;
      W_bmask_253_delayed_5_0_251_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_253_delayed_5_0_251_inst_req_1;
      W_bmask_253_delayed_5_0_251_inst_ack_1<= rack(0);
      W_bmask_253_delayed_5_0_251_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_253_delayed_5_0_251_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_253_delayed_5_0_253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_256_delayed_5_0_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_256_delayed_5_0_257_inst_req_0;
      W_index_256_delayed_5_0_257_inst_ack_0<= wack(0);
      rreq(0) <= W_index_256_delayed_5_0_257_inst_req_1;
      W_index_256_delayed_5_0_257_inst_ack_1<= rack(0);
      W_index_256_delayed_5_0_257_inst : InterlockBuffer generic map ( -- 
        name => "W_index_256_delayed_5_0_257_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_256_delayed_5_0_259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_252_delayed_5_0_248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_252_delayed_5_0_248_inst_req_0;
      W_rwbar_252_delayed_5_0_248_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_252_delayed_5_0_248_inst_req_1;
      W_rwbar_252_delayed_5_0_248_inst_ack_1<= rack(0);
      W_rwbar_252_delayed_5_0_248_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_252_delayed_5_0_248_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_252_delayed_5_0_250,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_260_delayed_5_0_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_260_delayed_5_0_267_inst_req_0;
      W_rwbar_260_delayed_5_0_267_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_260_delayed_5_0_267_inst_req_1;
      W_rwbar_260_delayed_5_0_267_inst_ack_1<= rack(0);
      W_rwbar_260_delayed_5_0_267_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_260_delayed_5_0_267_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_260_delayed_5_0_269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_255_delayed_5_0_254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_255_delayed_5_0_254_inst_req_0;
      W_wdata_255_delayed_5_0_254_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_255_delayed_5_0_254_inst_req_1;
      W_wdata_255_delayed_5_0_254_inst_ack_1<= rack(0);
      W_wdata_255_delayed_5_0_254_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_255_delayed_5_0_254_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_255_delayed_5_0_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nI_201_190_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_201_190_buf_req_0;
      nI_201_190_buf_ack_0<= wack(0);
      rreq(0) <= nI_201_190_buf_req_1;
      nI_201_190_buf_ack_1<= rack(0);
      nI_201_190_buf : InterlockBuffer generic map ( -- 
        name => "nI_201_190_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 7,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_201_190_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_193_addr_0
    process(array_obj_ref_193_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_193_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_193_gather_scatter
    process(type_cast_195_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_195_wire_constant;
      ov(31 downto 0) := iv;
      array_obj_ref_193_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_193_index_0_rename
    process(R_I_192_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_192_resized;
      ov(5 downto 0) := iv;
      R_I_192_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_193_index_0_resize
    process(I_185) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_185;
      ov := iv(5 downto 0);
      R_I_192_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_193_index_offset
    process(R_I_192_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_192_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_193_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_193_root_address_inst
    process(array_obj_ref_193_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_193_root_address <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_243_addr_0
    process(array_obj_ref_243_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_243_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_243_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_243_gather_scatter
    process(array_obj_ref_243_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_243_data_0;
      ov(31 downto 0) := iv;
      rval_244 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_243_index_0_rename
    process(R_index_242_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_242_resized;
      ov(5 downto 0) := iv;
      R_index_242_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_243_index_0_resize
    process(index_236) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_236;
      ov(5 downto 0) := iv;
      R_index_242_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_243_index_offset
    process(R_index_242_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_242_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_243_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_243_root_address_inst
    process(array_obj_ref_243_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_243_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_243_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_219_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_287_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_219_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_219_branch_req_0,
          ack0 => do_while_stmt_219_branch_ack_0,
          ack1 => do_while_stmt_219_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_210_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u7_u1_213_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_210_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_210_branch_req_0,
          ack0 => if_stmt_210_branch_ack_0,
          ack1 => if_stmt_210_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u7_u7_200_inst
    process(I_185) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_185, konst_199_wire_constant, tmp_var);
      nI_201 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_281_inst
    process(type_cast_279_wire_constant, rdata_276) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_279_wire_constant, rdata_276, tmp_var);
      resp_282 <= tmp_var; --
    end process;
    -- binary operator EQ_u7_u1_205_inst
    process(I_185) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_185, konst_204_wire_constant, tmp_var);
      EQ_u7_u1_205_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u7_u1_213_inst
    process(I_185) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(I_185, konst_212_wire_constant, tmp_var);
      ULT_u7_u1_213_wire <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_243_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_243_load_0_req_0;
      array_obj_ref_243_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_243_load_0_req_1;
      array_obj_ref_243_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_243_word_address_0;
      array_obj_ref_243_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : array_obj_ref_193_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_193_store_0_req_0;
      array_obj_ref_193_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_193_store_0_req_1;
      array_obj_ref_193_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_193_word_address_0;
      data_in <= array_obj_ref_193_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(5 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(42 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_req_0;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_req_1;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_222_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_223 <= data_out(42 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0", data_width => 43,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_MAC_ENABLE_202_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_MAC_ENABLE_202_inst_req_0;
      WPIPE_MAC_ENABLE_202_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_MAC_ENABLE_202_inst_req_1;
      WPIPE_MAC_ENABLE_202_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= MUX_208_wire;
      MAC_ENABLE_write_0_gI: SplitGuardInterface generic map(name => "MAC_ENABLE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      MAC_ENABLE_write_0: OutputPortRevised -- 
        generic map ( name => "MAC_ENABLE", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => MAC_ENABLE_pipe_write_req(0),
          oack => MAC_ENABLE_pipe_write_ack(0),
          odata => MAC_ENABLE_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_req_0;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_req_1;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_283_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_282;
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_1_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_1: OutputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_266_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_266_call_req_0;
      call_stmt_266_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_266_call_req_1;
      call_stmt_266_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_252_delayed_5_0_250(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_253_delayed_5_0_253 & rval_244 & wdata_255_delayed_5_0_256 & index_256_delayed_5_0_259;
      wval_266 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end NicRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    FREE_Q : in std_logic_vector(35 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(35 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_2109_start: Boolean;
  signal ReceiveEngineDaemon_CP_2109_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(54 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1539_call_req_0 : boolean;
  signal call_stmt_1539_call_ack_0 : boolean;
  signal NOT_u1_u1_1569_inst_req_0 : boolean;
  signal call_stmt_1556_call_ack_1 : boolean;
  signal call_stmt_1556_call_req_1 : boolean;
  signal NOT_u1_u1_1559_inst_ack_1 : boolean;
  signal call_stmt_1556_call_req_0 : boolean;
  signal call_stmt_1556_call_ack_0 : boolean;
  signal call_stmt_1593_call_ack_0 : boolean;
  signal NOT_u1_u1_1569_inst_ack_0 : boolean;
  signal call_stmt_1527_call_req_1 : boolean;
  signal ADD_u32_u32_1598_inst_req_1 : boolean;
  signal call_stmt_1527_call_ack_1 : boolean;
  signal NOT_u1_u1_1559_inst_req_1 : boolean;
  signal call_stmt_1593_call_ack_1 : boolean;
  signal npkt_cnt_1608_1517_buf_req_1 : boolean;
  signal npkt_cnt_1608_1517_buf_ack_1 : boolean;
  signal call_stmt_1593_call_req_1 : boolean;
  signal NOT_u1_u1_1559_inst_ack_0 : boolean;
  signal W_pkt_cnt_1581_delayed_13_0_1581_inst_req_0 : boolean;
  signal ADD_u32_u32_1598_inst_ack_0 : boolean;
  signal if_stmt_1505_branch_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_ack_0 : boolean;
  signal ADD_u32_u32_1598_inst_req_0 : boolean;
  signal if_stmt_1505_branch_ack_1 : boolean;
  signal NOT_u1_u1_1559_inst_req_0 : boolean;
  signal npkt_cnt_1608_1517_buf_ack_0 : boolean;
  signal npkt_cnt_1608_1517_buf_req_0 : boolean;
  signal NOT_u1_u1_1569_inst_ack_1 : boolean;
  signal NOT_u1_u1_1569_inst_req_1 : boolean;
  signal call_stmt_1527_call_ack_0 : boolean;
  signal ADD_u32_u32_1598_inst_ack_1 : boolean;
  signal W_pkt_cnt_1581_delayed_13_0_1581_inst_ack_1 : boolean;
  signal call_stmt_1527_call_req_0 : boolean;
  signal W_pkt_cnt_1590_delayed_13_0_1600_inst_req_0 : boolean;
  signal W_pkt_cnt_1590_delayed_13_0_1600_inst_req_1 : boolean;
  signal W_pkt_cnt_1590_delayed_13_0_1600_inst_ack_0 : boolean;
  signal do_while_stmt_1513_branch_req_0 : boolean;
  signal W_pkt_cnt_1590_delayed_13_0_1600_inst_ack_1 : boolean;
  signal call_stmt_1539_call_ack_1 : boolean;
  signal call_stmt_1539_call_req_1 : boolean;
  signal phi_stmt_1515_ack_0 : boolean;
  signal phi_stmt_1515_req_1 : boolean;
  signal call_stmt_1593_call_req_0 : boolean;
  signal W_pkt_cnt_1581_delayed_13_0_1581_inst_req_1 : boolean;
  signal phi_stmt_1515_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_req_1 : boolean;
  signal if_stmt_1505_branch_ack_0 : boolean;
  signal W_pkt_cnt_1581_delayed_13_0_1581_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_ack_1 : boolean;
  signal call_stmt_1618_call_req_0 : boolean;
  signal call_stmt_1618_call_ack_0 : boolean;
  signal call_stmt_1618_call_req_1 : boolean;
  signal call_stmt_1618_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_ack_1 : boolean;
  signal call_stmt_1631_call_req_0 : boolean;
  signal call_stmt_1631_call_ack_0 : boolean;
  signal call_stmt_1631_call_req_1 : boolean;
  signal call_stmt_1631_call_ack_1 : boolean;
  signal do_while_stmt_1513_branch_ack_0 : boolean;
  signal do_while_stmt_1513_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_2109_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_2109_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_2109_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_2109_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_2109: Block -- control-path 
    signal ReceiveEngineDaemon_CP_2109_elements: BooleanArray(91 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_2109_elements(0) <= ReceiveEngineDaemon_CP_2109_start;
    ReceiveEngineDaemon_CP_2109_symbol <= ReceiveEngineDaemon_CP_2109_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_sample_start_
      -- CP-element group 0: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Sample/req
      -- CP-element group 0: 	 assign_stmt_1501/$entry
      -- CP-element group 0: 	 $entry
      -- 
    req_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_update_start_
      -- CP-element group 1: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Update/req
      -- CP-element group 1: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Update/$entry
      -- 
    ack_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(1)); -- 
    req_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	91 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_update_completed_
      -- CP-element group 2: 	 assign_stmt_1501/$exit
      -- CP-element group 2: 	 branch_block_stmt_1502/merge_stmt_1504__entry__
      -- CP-element group 2: 	 branch_block_stmt_1502/$entry
      -- CP-element group 2: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Update/ack
      -- CP-element group 2: 	 assign_stmt_1501/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1502/branch_block_stmt_1502__entry__
      -- CP-element group 2: 	 branch_block_stmt_1502/merge_stmt_1504_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1502/merge_stmt_1504__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1502/merge_stmt_1504__entry___PhiReq/$exit
      -- 
    ack_2128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1502/$exit
      -- CP-element group 3: 	 branch_block_stmt_1502/branch_block_stmt_1502__exit__
      -- CP-element group 3: 	 $exit
      -- 
    ReceiveEngineDaemon_CP_2109_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	90 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	91 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1502/do_while_stmt_1513__exit__
      -- CP-element group 4: 	 branch_block_stmt_1502/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_1502/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1502/disable_loopback_PhiReq/$exit
      -- 
    ReceiveEngineDaemon_CP_2109_elements(4) <= ReceiveEngineDaemon_CP_2109_elements(90);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	91 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	91 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1502/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1502/if_stmt_1505_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1502/if_stmt_1505_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1502/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1502/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1505_branch_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	91 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_1502/do_while_stmt_1513__entry__
      -- CP-element group 6: 	 branch_block_stmt_1502/if_stmt_1505__exit__
      -- CP-element group 6: 	 branch_block_stmt_1502/if_stmt_1505_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1502/if_stmt_1505_else_link/$exit
      -- 
    else_choice_transition_2205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1505_branch_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513__entry__
      -- CP-element group 7: 	 branch_block_stmt_1502/do_while_stmt_1513/$entry
      -- 
    ReceiveEngineDaemon_CP_2109_elements(7) <= ReceiveEngineDaemon_CP_2109_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	90 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513__exit__
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_back
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	88 
    -- CP-element group 10: 	89 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1502/do_while_stmt_1513/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_taken/$entry
      -- 
    ReceiveEngineDaemon_CP_2109_elements(10) <= ReceiveEngineDaemon_CP_2109_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	87 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_body_done
      -- 
    ReceiveEngineDaemon_CP_2109_elements(11) <= ReceiveEngineDaemon_CP_2109_elements(87);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/back_edge_to_loop_body
      -- 
    ReceiveEngineDaemon_CP_2109_elements(12) <= ReceiveEngineDaemon_CP_2109_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	23 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/first_time_through_loop_body
      -- 
    ReceiveEngineDaemon_CP_2109_elements(13) <= ReceiveEngineDaemon_CP_2109_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	34 
    -- CP-element group 14: 	86 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	18 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/$entry
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	86 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/condition_evaluated
      -- 
    condition_evaluated_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(15), ack => do_while_stmt_1513_branch_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(86) & ReceiveEngineDaemon_CP_2109_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_sample_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(17) & ReceiveEngineDaemon_CP_2109_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	65 
    -- CP-element group 17: 	69 
    -- CP-element group 17: 	45 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	16 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_sample_start_
      -- 
    ReceiveEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(14) & ReceiveEngineDaemon_CP_2109_elements(65) & ReceiveEngineDaemon_CP_2109_elements(69) & ReceiveEngineDaemon_CP_2109_elements(45) & ReceiveEngineDaemon_CP_2109_elements(49) & ReceiveEngineDaemon_CP_2109_elements(19);
      gj_ReceiveEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	68 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_update_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(14) & ReceiveEngineDaemon_CP_2109_elements(56) & ReceiveEngineDaemon_CP_2109_elements(64) & ReceiveEngineDaemon_CP_2109_elements(68);
      gj_ReceiveEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	67 
    -- CP-element group 19: 	43 
    -- CP-element group 19: 	47 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_sample_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	54 
    -- CP-element group 20: 	62 
    -- CP-element group 20: 	66 
    -- CP-element group 20: 	15 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/aggregated_phi_update_ack
      -- CP-element group 20: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_update_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	12 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_loopback_trigger
      -- 
    ReceiveEngineDaemon_CP_2109_elements(21) <= ReceiveEngineDaemon_CP_2109_elements(12);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_loopback_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_loopback_sample_req
      -- 
    phi_stmt_1515_loopback_sample_req_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_loopback_sample_req_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(22), ack => phi_stmt_1515_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	13 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_entry_trigger
      -- 
    ReceiveEngineDaemon_CP_2109_elements(23) <= ReceiveEngineDaemon_CP_2109_elements(13);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_entry_sample_req
      -- 
    phi_stmt_1515_entry_sample_req_2239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_entry_sample_req_2239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(24), ack => phi_stmt_1515_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_phi_mux_ack_ps
      -- CP-element group 25: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/phi_stmt_1515_phi_mux_ack
      -- 
    phi_stmt_1515_phi_mux_ack_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1515_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Sample/req
      -- CP-element group 26: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_sample_start__ps
      -- 
    req_2255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(26), ack => npkt_cnt_1608_1517_buf_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Update/req
      -- CP-element group 27: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_update_start__ps
      -- 
    req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(27), ack => npkt_cnt_1608_1517_buf_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_sample_completed__ps
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1608_1517_buf_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Update/ack
      -- CP-element group 29: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/R_npkt_cnt_1517_update_completed__ps
      -- 
    ack_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1608_1517_buf_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_sample_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_update_start_
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_update_completed__ps
      -- 
    ReceiveEngineDaemon_CP_2109_elements(32) <= ReceiveEngineDaemon_CP_2109_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/type_cast_1519_update_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_2109_elements(31), ack => ReceiveEngineDaemon_CP_2109_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	14 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	85 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Sample/crr
      -- CP-element group 34: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_sample_start_
      -- 
    crr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(34), ack => call_stmt_1527_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(14) & ReceiveEngineDaemon_CP_2109_elements(36) & ReceiveEngineDaemon_CP_2109_elements(85);
      gj_ReceiveEngineDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	52 
    -- CP-element group 35: 	72 
    -- CP-element group 35: 	80 
    -- CP-element group 35: 	85 
    -- CP-element group 35: 	40 
    -- CP-element group 35: 	44 
    -- CP-element group 35: 	48 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Update/ccr
      -- CP-element group 35: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_update_start_
      -- 
    ccr_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(35), ack => call_stmt_1527_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(52) & ReceiveEngineDaemon_CP_2109_elements(72) & ReceiveEngineDaemon_CP_2109_elements(80) & ReceiveEngineDaemon_CP_2109_elements(85) & ReceiveEngineDaemon_CP_2109_elements(40) & ReceiveEngineDaemon_CP_2109_elements(44) & ReceiveEngineDaemon_CP_2109_elements(48);
      gj_ReceiveEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Sample/cra
      -- CP-element group 36: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_sample_completed_
      -- 
    cra_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1527_call_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	42 
    -- CP-element group 37: 	46 
    -- CP-element group 37: 	50 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1527_update_completed_
      -- 
    cca_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1527_call_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	77 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Sample/crr
      -- CP-element group 38: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_sample_start_
      -- 
    crr_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(38), ack => call_stmt_1539_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(37) & ReceiveEngineDaemon_CP_2109_elements(77) & ReceiveEngineDaemon_CP_2109_elements(40);
      gj_ReceiveEngineDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	77 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Update/ccr
      -- 
    ccr_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(39), ack => call_stmt_1539_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(77) & ReceiveEngineDaemon_CP_2109_elements(41);
      gj_ReceiveEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	35 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Sample/cra
      -- CP-element group 40: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_sample_completed_
      -- 
    cra_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1539_call_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Update/cca
      -- CP-element group 41: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1539_Update/$exit
      -- 
    cca_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1539_call_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Sample/crr
      -- CP-element group 42: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_sample_start_
      -- 
    crr_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(42), ack => call_stmt_1556_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(37) & ReceiveEngineDaemon_CP_2109_elements(44);
      gj_ReceiveEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	19 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	60 
    -- CP-element group 43: 	76 
    -- CP-element group 43: 	84 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Update/ccr
      -- CP-element group 43: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_update_start_
      -- 
    ccr_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(43), ack => call_stmt_1556_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(19) & ReceiveEngineDaemon_CP_2109_elements(60) & ReceiveEngineDaemon_CP_2109_elements(76) & ReceiveEngineDaemon_CP_2109_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Sample/cra
      -- CP-element group 44: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_sample_completed_
      -- 
    cra_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1556_call_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45: 	74 
    -- CP-element group 45: 	82 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	17 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Update/cca
      -- CP-element group 45: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1556_update_completed_
      -- 
    cca_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1556_call_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	37 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Sample/$entry
      -- 
    rr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(46), ack => NOT_u1_u1_1559_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(37) & ReceiveEngineDaemon_CP_2109_elements(48);
      gj_ReceiveEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	19 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	60 
    -- CP-element group 47: 	76 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Update/cr
      -- CP-element group 47: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_update_start_
      -- 
    cr_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(47), ack => NOT_u1_u1_1559_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(19) & ReceiveEngineDaemon_CP_2109_elements(60) & ReceiveEngineDaemon_CP_2109_elements(76);
      gj_ReceiveEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Sample/$exit
      -- 
    ra_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1559_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49: 	74 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	17 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1559_update_completed_
      -- 
    ca_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1559_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	37 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_sample_start_
      -- 
    rr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(50), ack => NOT_u1_u1_1569_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(37) & ReceiveEngineDaemon_CP_2109_elements(52);
      gj_ReceiveEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	84 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Update/cr
      -- 
    cr_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(51), ack => NOT_u1_u1_1569_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	35 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_sample_completed_
      -- 
    ra_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1569_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	82 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/NOT_u1_u1_1569_Update/ca
      -- 
    ca_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1569_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	20 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Sample/req
      -- 
    req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(54), ack => W_pkt_cnt_1581_delayed_13_0_1581_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(20) & ReceiveEngineDaemon_CP_2109_elements(56);
      gj_ReceiveEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Update/req
      -- CP-element group 55: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Update/$entry
      -- 
    req_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(55), ack => W_pkt_cnt_1581_delayed_13_0_1581_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	18 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Sample/ack
      -- 
    ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1581_delayed_13_0_1581_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Update/ack
      -- CP-element group 57: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1583_Update/$exit
      -- 
    ack_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1581_delayed_13_0_1581_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	49 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Sample/crr
      -- 
    crr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(58), ack => call_stmt_1593_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 31,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(57) & ReceiveEngineDaemon_CP_2109_elements(41) & ReceiveEngineDaemon_CP_2109_elements(45) & ReceiveEngineDaemon_CP_2109_elements(49) & ReceiveEngineDaemon_CP_2109_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_update_start_
      -- 
    ccr_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(59), ack => call_stmt_1593_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(61);
      gj_ReceiveEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	43 
    -- CP-element group 60: 	47 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Sample/cra
      -- CP-element group 60: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_sample_completed_
      -- 
    cra_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1593_call_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	74 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Update/cca
      -- CP-element group 61: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1593_update_completed_
      -- 
    cca_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1593_call_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	20 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Sample/$entry
      -- 
    rr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(62), ack => ADD_u32_u32_1598_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(20) & ReceiveEngineDaemon_CP_2109_elements(64);
      gj_ReceiveEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Update/$entry
      -- 
    cr_2381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(63), ack => ADD_u32_u32_1598_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(19) & ReceiveEngineDaemon_CP_2109_elements(65);
      gj_ReceiveEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	18 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Sample/ra
      -- CP-element group 64: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Sample/$exit
      -- 
    ra_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1598_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	87 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	17 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/ADD_u32_u32_1598_update_completed_
      -- 
    ca_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1598_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	20 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Sample/req
      -- CP-element group 66: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_sample_start_
      -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(66), ack => W_pkt_cnt_1590_delayed_13_0_1600_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(20) & ReceiveEngineDaemon_CP_2109_elements(68);
      gj_ReceiveEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	19 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Update/req
      -- CP-element group 67: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_update_start_
      -- 
    req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(67), ack => W_pkt_cnt_1590_delayed_13_0_1600_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(19) & ReceiveEngineDaemon_CP_2109_elements(69);
      gj_ReceiveEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	18 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Sample/$exit
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1590_delayed_13_0_1600_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	87 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	17 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1602_Update/ack
      -- 
    ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1590_delayed_13_0_1600_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Sample/req
      -- 
    req_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(70), ack => W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(37) & ReceiveEngineDaemon_CP_2109_elements(72);
      gj_ReceiveEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	76 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Update/req
      -- 
    req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(71), ack => W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(76);
      gj_ReceiveEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	35 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Sample/ack
      -- 
    ack_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1615_Update/ack
      -- 
    ack_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	61 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	45 
    -- CP-element group 74: 	49 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Sample/crr
      -- 
    crr_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(74), ack => call_stmt_1618_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(61) & ReceiveEngineDaemon_CP_2109_elements(73) & ReceiveEngineDaemon_CP_2109_elements(45) & ReceiveEngineDaemon_CP_2109_elements(49) & ReceiveEngineDaemon_CP_2109_elements(76);
      gj_ReceiveEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Update/ccr
      -- 
    ccr_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(75), ack => call_stmt_1618_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(77);
      gj_ReceiveEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	43 
    -- CP-element group 76: 	47 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Sample/cra
      -- 
    cra_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1618_call_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	38 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	39 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1618_Update/cca
      -- 
    cca_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1618_call_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Sample/req
      -- 
    req_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(78), ack => W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(37) & ReceiveEngineDaemon_CP_2109_elements(80);
      gj_ReceiveEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	84 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_update_start_
      -- CP-element group 79: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Update/req
      -- 
    req_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(79), ack => W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	35 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Sample/ack
      -- 
    ack_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/assign_stmt_1623_Update/ack
      -- 
    ack_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	53 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	81 
    -- CP-element group 82: 	45 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Sample/crr
      -- 
    crr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(82), ack => call_stmt_1631_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 31,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(53) & ReceiveEngineDaemon_CP_2109_elements(77) & ReceiveEngineDaemon_CP_2109_elements(81) & ReceiveEngineDaemon_CP_2109_elements(45) & ReceiveEngineDaemon_CP_2109_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_update_start_
      -- CP-element group 83: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Update/ccr
      -- 
    ccr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(83), ack => call_stmt_1631_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2109_elements(85);
      gj_ReceiveEngineDaemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	51 
    -- CP-element group 84: 	79 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	43 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Sample/cra
      -- 
    cra_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1631_call_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	34 
    -- CP-element group 85: 	35 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/call_stmt_1631_Update/cca
      -- 
    cca_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1631_call_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	14 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	15 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_2109_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_2109_elements(14), ack => ReceiveEngineDaemon_CP_2109_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	65 
    -- CP-element group 87: 	69 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	11 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1502/do_while_stmt_1513/do_while_stmt_1513_loop_body/$exit
      -- 
    ReceiveEngineDaemon_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2109_elements(65) & ReceiveEngineDaemon_CP_2109_elements(69) & ReceiveEngineDaemon_CP_2109_elements(85);
      gj_ReceiveEngineDaemon_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	10 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_exit/$exit
      -- CP-element group 88: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_exit/ack
      -- 
    ack_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1513_branch_ack_0, ack => ReceiveEngineDaemon_CP_2109_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	10 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_taken/$exit
      -- CP-element group 89: 	 branch_block_stmt_1502/do_while_stmt_1513/loop_taken/ack
      -- 
    ack_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1513_branch_ack_1, ack => ReceiveEngineDaemon_CP_2109_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	8 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	4 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1502/do_while_stmt_1513/$exit
      -- 
    ReceiveEngineDaemon_CP_2109_elements(90) <= ReceiveEngineDaemon_CP_2109_elements(8);
    -- CP-element group 91:  merge  branch  transition  place  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	2 
    -- CP-element group 91: 	4 
    -- CP-element group 91: 	5 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	5 
    -- CP-element group 91: 	6 
    -- CP-element group 91:  members (49) 
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Update/ack
      -- CP-element group 91: 	 branch_block_stmt_1502/NOT_u1_u1_1509_place
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Update/cr
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Update/req
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Sample/req
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/branch_req
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_if_link/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/SplitProtocol/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Update/cr
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/BITSEL_u32_u1_1508_inputs/RPIPE_CONTROL_REGISTER_1506/Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505__entry__
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_eval_test/NOT_u1_u1_1509/BITSEL_u32_u1_1508/SplitProtocol/Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/merge_stmt_1504__exit__
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_dead_link/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/if_stmt_1505_else_link/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/merge_stmt_1504_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_1502/merge_stmt_1504_PhiAck/$entry
      -- CP-element group 91: 	 branch_block_stmt_1502/merge_stmt_1504_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_1502/merge_stmt_1504_PhiAck/dummy
      -- 
    branch_req_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2109_elements(91), ack => if_stmt_1505_branch_req_0); -- 
    ReceiveEngineDaemon_CP_2109_elements(91) <= OrReduce(ReceiveEngineDaemon_CP_2109_elements(2) & ReceiveEngineDaemon_CP_2109_elements(4) & ReceiveEngineDaemon_CP_2109_elements(5));
    ReceiveEngineDaemon_do_while_stmt_1513_terminator_2462: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_1513_terminator_2462", max_iterations_in_flight =>31) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_2109_elements(11),loop_continue => ReceiveEngineDaemon_CP_2109_elements(89),loop_terminate => ReceiveEngineDaemon_CP_2109_elements(88),loop_back => ReceiveEngineDaemon_CP_2109_elements(9),loop_exit => ReceiveEngineDaemon_CP_2109_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1515_phi_seq_2270_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ReceiveEngineDaemon_CP_2109_elements(21);
      ReceiveEngineDaemon_CP_2109_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ReceiveEngineDaemon_CP_2109_elements(28);
      ReceiveEngineDaemon_CP_2109_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= ReceiveEngineDaemon_CP_2109_elements(29);
      ReceiveEngineDaemon_CP_2109_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= ReceiveEngineDaemon_CP_2109_elements(23);
      ReceiveEngineDaemon_CP_2109_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ReceiveEngineDaemon_CP_2109_elements(30);
      ReceiveEngineDaemon_CP_2109_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= ReceiveEngineDaemon_CP_2109_elements(32);
      ReceiveEngineDaemon_CP_2109_elements(24) <= phi_mux_reqs(1);
      phi_stmt_1515_phi_seq_2270 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1515_phi_seq_2270") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ReceiveEngineDaemon_CP_2109_elements(16), 
          phi_sample_ack => ReceiveEngineDaemon_CP_2109_elements(19), 
          phi_update_req => ReceiveEngineDaemon_CP_2109_elements(18), 
          phi_update_ack => ReceiveEngineDaemon_CP_2109_elements(20), 
          phi_mux_ack => ReceiveEngineDaemon_CP_2109_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2222_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_2109_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_2109_elements(13);
        entry_tmerge_2222 : transition_merge -- 
          generic map(name => " entry_tmerge_2222")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_2109_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1589_1589_delayed_13_0_1599 : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_1508_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1636_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1509_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1558_1558_delayed_10_0_1560 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1564_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1565_1565_delayed_10_0_1570 : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1535_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1589_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1506_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1634_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1524_wire : std_logic_vector(35 downto 0);
    signal RPIPE_FREE_Q_1627_wire : std_logic_vector(35 downto 0);
    signal bad_packet_identifier_1556 : std_logic_vector(0 downto 0);
    signal cond_1580 : std_logic_vector(0 downto 0);
    signal free_flag_1575 : std_logic_vector(0 downto 0);
    signal ignore_resp0_1539 : std_logic_vector(31 downto 0);
    signal ignore_resp1_1593 : std_logic_vector(31 downto 0);
    signal konst_1500_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1507_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1536_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1578_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1590_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1635_wire_constant : std_logic_vector(31 downto 0);
    signal npkt_cnt_1608 : std_logic_vector(31 downto 0);
    signal npkt_cnt_1608_1517_buffered : std_logic_vector(31 downto 0);
    signal ok_flag_1566 : std_logic_vector(0 downto 0);
    signal pkt_cnt_1515 : std_logic_vector(31 downto 0);
    signal pkt_cnt_1581_delayed_13_0_1583 : std_logic_vector(31 downto 0);
    signal pkt_cnt_1590_delayed_13_0_1602 : std_logic_vector(31 downto 0);
    signal push_status_1631 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_32_1527 : std_logic_vector(31 downto 0);
    signal rx_buffer_pointer_36_1545 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1598_delayed_10_0_1615 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1606_delayed_10_0_1623 : std_logic_vector(35 downto 0);
    signal slice_1629_wire : std_logic_vector(31 downto 0);
    signal status_1527 : std_logic_vector(0 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1523_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1532_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1542_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1586_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1626_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1535_wire_constant <= "1111";
    NOT_u4_u4_1589_wire_constant <= "1111";
    konst_1500_wire_constant <= "000000";
    konst_1507_wire_constant <= "00000000000000000000000000000000";
    konst_1536_wire_constant <= "011000";
    konst_1578_wire_constant <= "1";
    konst_1590_wire_constant <= "011001";
    konst_1635_wire_constant <= "00000000000000000000000000000000";
    type_cast_1519_wire_constant <= "00000000000000000000000000000000";
    type_cast_1523_wire_constant <= "1";
    type_cast_1532_wire_constant <= "0";
    type_cast_1542_wire_constant <= "0000";
    type_cast_1586_wire_constant <= "0";
    type_cast_1597_wire_constant <= "00000000000000000000000000000001";
    type_cast_1626_wire_constant <= "1";
    phi_stmt_1515: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= npkt_cnt_1608_1517_buffered & type_cast_1519_wire_constant;
      req <= phi_stmt_1515_req_0 & phi_stmt_1515_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1515",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1515_ack_0,
          idata => idata,
          odata => pkt_cnt_1515,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1515
    -- flow-through select operator MUX_1607_inst
    npkt_cnt_1608 <= ADD_u32_u32_1589_1589_delayed_13_0_1599 when (ok_flag_1566(0) /=  '0') else pkt_cnt_1590_delayed_13_0_1602;
    -- flow-through slice operator slice_1629_inst
    slice_1629_wire <= rx_buffer_pointer_36_1606_delayed_10_0_1623(31 downto 0);
    W_pkt_cnt_1581_delayed_13_0_1581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_cnt_1581_delayed_13_0_1581_inst_req_0;
      W_pkt_cnt_1581_delayed_13_0_1581_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_cnt_1581_delayed_13_0_1581_inst_req_1;
      W_pkt_cnt_1581_delayed_13_0_1581_inst_ack_1<= rack(0);
      W_pkt_cnt_1581_delayed_13_0_1581_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_cnt_1581_delayed_13_0_1581_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_cnt_1515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_cnt_1581_delayed_13_0_1583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_cnt_1590_delayed_13_0_1600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_cnt_1590_delayed_13_0_1600_inst_req_0;
      W_pkt_cnt_1590_delayed_13_0_1600_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_cnt_1590_delayed_13_0_1600_inst_req_1;
      W_pkt_cnt_1590_delayed_13_0_1600_inst_ack_1<= rack(0);
      W_pkt_cnt_1590_delayed_13_0_1600_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_cnt_1590_delayed_13_0_1600_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_cnt_1515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_cnt_1590_delayed_13_0_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_req_0;
      W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_req_1;
      W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1598_delayed_10_0_1613_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_1545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1598_delayed_10_0_1615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_req_0;
      W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_req_1;
      W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1606_delayed_10_0_1621_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_1545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1606_delayed_10_0_1623,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_1608_1517_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_1608_1517_buf_req_0;
      npkt_cnt_1608_1517_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_1608_1517_buf_req_1;
      npkt_cnt_1608_1517_buf_ack_1<= rack(0);
      npkt_cnt_1608_1517_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_1608_1517_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_1608_1517_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1513_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1636_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1513_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1513_branch_req_0,
          ack0 => do_while_stmt_1513_branch_ack_0,
          ack1 => do_while_stmt_1513_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1505_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1509_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1505_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1505_branch_req_0,
          ack0 => if_stmt_1505_branch_ack_0,
          ack1 => if_stmt_1505_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_1598_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 13);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pkt_cnt_1515;
      ADD_u32_u32_1589_1589_delayed_13_0_1599 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_1598_inst_req_0;
      ADD_u32_u32_1598_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_1598_inst_req_1;
      ADD_u32_u32_1598_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 13,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator AND_u1_u1_1565_inst
    process(NOT_u1_u1_1558_1558_delayed_10_0_1560, NOT_u1_u1_1564_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1558_1558_delayed_10_0_1560, NOT_u1_u1_1564_wire, tmp_var);
      ok_flag_1566 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1574_inst
    process(NOT_u1_u1_1565_1565_delayed_10_0_1570, bad_packet_identifier_1556) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1565_1565_delayed_10_0_1570, bad_packet_identifier_1556, tmp_var);
      free_flag_1575 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1508_inst
    process(RPIPE_CONTROL_REGISTER_1506_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1506_wire, konst_1507_wire_constant, tmp_var);
      BITSEL_u32_u1_1508_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1636_inst
    process(RPIPE_CONTROL_REGISTER_1634_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1634_wire, konst_1635_wire_constant, tmp_var);
      BITSEL_u32_u1_1636_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1544_inst
    process(type_cast_1542_wire_constant, rx_buffer_pointer_32_1527) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1542_wire_constant, rx_buffer_pointer_32_1527, tmp_var);
      rx_buffer_pointer_36_1545 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1579_inst
    process(ok_flag_1566) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ok_flag_1566, konst_1578_wire_constant, tmp_var);
      cond_1580 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1509_inst
    process(BITSEL_u32_u1_1508_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1508_wire, tmp_var);
      NOT_u1_u1_1509_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (8) : NOT_u1_u1_1559_inst 
    ApIntNot_group_8: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1527;
      NOT_u1_u1_1558_1558_delayed_10_0_1560 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1559_inst_req_0;
      NOT_u1_u1_1559_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1559_inst_req_1;
      NOT_u1_u1_1559_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_8_gI: SplitGuardInterface generic map(name => "ApIntNot_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- unary operator NOT_u1_u1_1564_inst
    process(bad_packet_identifier_1556) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_1556, tmp_var);
      NOT_u1_u1_1564_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (10) : NOT_u1_u1_1569_inst 
    ApIntNot_group_10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1527;
      NOT_u1_u1_1565_1565_delayed_10_0_1570 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1569_inst_req_0;
      NOT_u1_u1_1569_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1569_inst_req_1;
      NOT_u1_u1_1569_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_10_gI: SplitGuardInterface generic map(name => "ApIntNot_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1506_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1634_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1524_wire <= FREE_Q;
    RPIPE_FREE_Q_1627_wire <= FREE_Q;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1499_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1500_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1527_call 
    popFromQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1527_call_req_0;
      call_stmt_1527_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1527_call_req_1;
      call_stmt_1527_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_0_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1523_wire_constant & RPIPE_FREE_Q_1524_wire;
      rx_buffer_pointer_32_1527 <= data_out(32 downto 1);
      status_1527 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1539_call call_stmt_1593_call 
    AccessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 4);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1539_call_req_0;
      reqL_unguarded(0) <= call_stmt_1593_call_req_0;
      call_stmt_1539_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1593_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1539_call_req_1;
      reqR_unguarded(0) <= call_stmt_1593_call_req_1;
      call_stmt_1539_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1593_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1566(0);
      guard_vector(1)  <=  not status_1527(0);
      AccessRegister_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1532_wire_constant & NOT_u4_u4_1535_wire_constant & konst_1536_wire_constant & rx_buffer_pointer_32_1527 & type_cast_1586_wire_constant & NOT_u4_u4_1589_wire_constant & konst_1590_wire_constant & pkt_cnt_1581_delayed_13_0_1583;
      ignore_resp0_1539 <= data_out(63 downto 32);
      ignore_resp1_1593 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1556_call 
    loadBuffer_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1556_call_req_0;
      call_stmt_1556_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1556_call_req_1;
      call_stmt_1556_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_1527(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_2_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1545;
      bad_packet_identifier_1556 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(35 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1618_call 
    populateRxQueue_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1618_call_req_0;
      call_stmt_1618_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1618_call_req_1;
      call_stmt_1618_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1566(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_3_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1598_delayed_10_0_1615;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(35 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1631_call 
    pushIntoQueue_call_group_4: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1631_call_req_0;
      call_stmt_1631_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1631_call_req_1;
      call_stmt_1631_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_1575(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_4_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1626_wire_constant & RPIPE_FREE_Q_1627_wire & slice_1629_wire;
      push_status_1631 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity SoftwareRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    MAC_ENABLE : in std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    enable_mac_pipe_write_req : out  std_logic_vector(0 downto 0);
    enable_mac_pipe_write_ack : in   std_logic_vector(0 downto 0);
    enable_mac_pipe_write_data : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity SoftwareRegisterAccessDaemon;
architecture SoftwareRegisterAccessDaemon_arch of SoftwareRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal SoftwareRegisterAccessDaemon_CP_2481_start: Boolean;
  signal SoftwareRegisterAccessDaemon_CP_2481_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal check_free_q_1783_1669_buf_ack_1 : boolean;
  signal check_control_regsiter_1774_1664_buf_req_0 : boolean;
  signal phi_stmt_1670_req_1 : boolean;
  signal check_control_regsiter_1774_1664_buf_req_1 : boolean;
  signal check_num_server_1792_1674_buf_req_1 : boolean;
  signal check_free_q_1783_1669_buf_req_1 : boolean;
  signal if_stmt_1646_branch_ack_0 : boolean;
  signal check_control_regsiter_1774_1664_buf_ack_1 : boolean;
  signal if_stmt_1646_branch_ack_1 : boolean;
  signal check_free_q_1783_1669_buf_ack_0 : boolean;
  signal check_free_q_1783_1669_buf_req_0 : boolean;
  signal check_num_server_1792_1674_buf_req_0 : boolean;
  signal phi_stmt_1660_req_1 : boolean;
  signal check_control_regsiter_1774_1664_buf_ack_0 : boolean;
  signal phi_stmt_1670_ack_0 : boolean;
  signal phi_stmt_1665_ack_0 : boolean;
  signal phi_stmt_1654_req_0 : boolean;
  signal phi_stmt_1654_req_1 : boolean;
  signal phi_stmt_1654_ack_0 : boolean;
  signal array_obj_ref_1710_load_0_req_0 : boolean;
  signal phi_stmt_1665_req_0 : boolean;
  signal phi_stmt_1670_req_0 : boolean;
  signal do_while_stmt_1652_branch_req_0 : boolean;
  signal check_num_server_1792_1674_buf_ack_0 : boolean;
  signal if_stmt_1646_branch_req_0 : boolean;
  signal array_obj_ref_1679_load_0_ack_0 : boolean;
  signal check_num_server_1792_1674_buf_ack_1 : boolean;
  signal phi_stmt_1660_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1708_inst_ack_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1708_inst_req_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1708_inst_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1708_inst_ack_0 : boolean;
  signal array_obj_ref_1679_load_0_ack_1 : boolean;
  signal array_obj_ref_1679_load_0_req_1 : boolean;
  signal array_obj_ref_1679_load_0_req_0 : boolean;
  signal array_obj_ref_1710_load_0_ack_1 : boolean;
  signal W_update_control_register_pipe_1690_delayed_5_0_1712_inst_req_0 : boolean;
  signal W_update_control_register_pipe_1690_delayed_5_0_1712_inst_ack_0 : boolean;
  signal array_obj_ref_1710_load_0_ack_0 : boolean;
  signal phi_stmt_1665_req_1 : boolean;
  signal phi_stmt_1660_req_0 : boolean;
  signal W_update_control_register_pipe_1690_delayed_5_0_1712_inst_req_1 : boolean;
  signal W_update_control_register_pipe_1690_delayed_5_0_1712_inst_ack_1 : boolean;
  signal array_obj_ref_1710_load_0_req_1 : boolean;
  signal array_obj_ref_1718_load_0_req_0 : boolean;
  signal array_obj_ref_1718_load_0_ack_0 : boolean;
  signal array_obj_ref_1718_load_0_req_1 : boolean;
  signal array_obj_ref_1718_load_0_ack_1 : boolean;
  signal EQ_u32_u1_1721_inst_req_0 : boolean;
  signal EQ_u32_u1_1721_inst_ack_0 : boolean;
  signal EQ_u32_u1_1721_inst_req_1 : boolean;
  signal EQ_u32_u1_1721_inst_ack_1 : boolean;
  signal WPIPE_enable_mac_1716_inst_req_0 : boolean;
  signal WPIPE_enable_mac_1716_inst_ack_0 : boolean;
  signal WPIPE_enable_mac_1716_inst_req_1 : boolean;
  signal WPIPE_enable_mac_1716_inst_ack_1 : boolean;
  signal array_obj_ref_1726_load_0_req_0 : boolean;
  signal array_obj_ref_1726_load_0_ack_0 : boolean;
  signal array_obj_ref_1726_load_0_req_1 : boolean;
  signal array_obj_ref_1726_load_0_ack_1 : boolean;
  signal W_update_free_q_pipe_1703_delayed_5_0_1728_inst_req_0 : boolean;
  signal W_update_free_q_pipe_1703_delayed_5_0_1728_inst_ack_0 : boolean;
  signal W_update_free_q_pipe_1703_delayed_5_0_1728_inst_req_1 : boolean;
  signal W_update_free_q_pipe_1703_delayed_5_0_1728_inst_ack_1 : boolean;
  signal type_cast_1734_inst_req_0 : boolean;
  signal type_cast_1734_inst_ack_0 : boolean;
  signal type_cast_1734_inst_req_1 : boolean;
  signal type_cast_1734_inst_ack_1 : boolean;
  signal WPIPE_FREE_Q_1732_inst_req_0 : boolean;
  signal WPIPE_FREE_Q_1732_inst_ack_0 : boolean;
  signal WPIPE_FREE_Q_1732_inst_req_1 : boolean;
  signal WPIPE_FREE_Q_1732_inst_ack_1 : boolean;
  signal array_obj_ref_1739_load_0_req_0 : boolean;
  signal array_obj_ref_1739_load_0_ack_0 : boolean;
  signal array_obj_ref_1739_load_0_req_1 : boolean;
  signal array_obj_ref_1739_load_0_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1737_inst_req_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1737_inst_ack_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1737_inst_req_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1737_inst_ack_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1742_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1742_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1742_inst_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1742_inst_ack_1 : boolean;
  signal array_obj_ref_1795_load_0_req_0 : boolean;
  signal array_obj_ref_1795_load_0_ack_0 : boolean;
  signal array_obj_ref_1795_load_0_req_1 : boolean;
  signal array_obj_ref_1795_load_0_ack_1 : boolean;
  signal W_index_1777_delayed_5_0_1797_inst_req_0 : boolean;
  signal W_index_1777_delayed_5_0_1797_inst_ack_0 : boolean;
  signal W_index_1777_delayed_5_0_1797_inst_req_1 : boolean;
  signal W_index_1777_delayed_5_0_1797_inst_ack_1 : boolean;
  signal W_wdata_1776_delayed_5_0_1800_inst_req_0 : boolean;
  signal W_wdata_1776_delayed_5_0_1800_inst_ack_0 : boolean;
  signal W_wdata_1776_delayed_5_0_1800_inst_req_1 : boolean;
  signal W_wdata_1776_delayed_5_0_1800_inst_ack_1 : boolean;
  signal W_bmask_1774_delayed_5_0_1803_inst_req_0 : boolean;
  signal W_bmask_1774_delayed_5_0_1803_inst_ack_0 : boolean;
  signal W_bmask_1774_delayed_5_0_1803_inst_req_1 : boolean;
  signal W_bmask_1774_delayed_5_0_1803_inst_ack_1 : boolean;
  signal W_rwbar_1773_delayed_5_0_1806_inst_req_0 : boolean;
  signal W_rwbar_1773_delayed_5_0_1806_inst_ack_0 : boolean;
  signal W_rwbar_1773_delayed_5_0_1806_inst_req_1 : boolean;
  signal W_rwbar_1773_delayed_5_0_1806_inst_ack_1 : boolean;
  signal call_stmt_1815_call_req_0 : boolean;
  signal call_stmt_1815_call_ack_0 : boolean;
  signal call_stmt_1815_call_req_1 : boolean;
  signal call_stmt_1815_call_ack_1 : boolean;
  signal W_rwbar_1781_delayed_5_0_1816_inst_req_0 : boolean;
  signal W_rwbar_1781_delayed_5_0_1816_inst_ack_0 : boolean;
  signal W_rwbar_1781_delayed_5_0_1816_inst_req_1 : boolean;
  signal W_rwbar_1781_delayed_5_0_1816_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1832_inst_req_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1832_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1832_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1832_inst_ack_1 : boolean;
  signal do_while_stmt_1652_branch_ack_0 : boolean;
  signal do_while_stmt_1652_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  SoftwareRegisterAccessDaemon_CP_2481_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2481_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2481_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2481_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  SoftwareRegisterAccessDaemon_CP_2481: Block -- control-path 
    signal SoftwareRegisterAccessDaemon_CP_2481_elements: BooleanArray(185 downto 0);
    -- 
  begin -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(0) <= SoftwareRegisterAccessDaemon_CP_2481_start;
    SoftwareRegisterAccessDaemon_CP_2481_symbol <= SoftwareRegisterAccessDaemon_CP_2481_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	185 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1642/merge_stmt_1643__entry__
      -- CP-element group 0: 	 branch_block_stmt_1642/branch_block_stmt_1642__entry__
      -- CP-element group 0: 	 branch_block_stmt_1642/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1642/merge_stmt_1643_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1642/merge_stmt_1643__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1642/merge_stmt_1643__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	184 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1642/do_while_stmt_1652__exit__
      -- CP-element group 1: 	 branch_block_stmt_1642/branch_block_stmt_1642__exit__
      -- CP-element group 1: 	 branch_block_stmt_1642/$exit
      -- CP-element group 1: 	 $exit
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(184);
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	185 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	185 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_1642/if_stmt_1646_if_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_1642/if_stmt_1646_if_link/if_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_1642/not_mac_enable_loopback
      -- CP-element group 2: 	 branch_block_stmt_1642/not_mac_enable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1642/not_mac_enable_loopback_PhiReq/$exit
      -- 
    if_choice_transition_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1646_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(2)); -- 
    -- CP-element group 3:  merge  transition  place  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	185 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (4) 
      -- CP-element group 3: 	 branch_block_stmt_1642/if_stmt_1646_else_link/else_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_1642/do_while_stmt_1652__entry__
      -- CP-element group 3: 	 branch_block_stmt_1642/if_stmt_1646__exit__
      -- CP-element group 3: 	 branch_block_stmt_1642/if_stmt_1646_else_link/$exit
      -- 
    else_choice_transition_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1646_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(3)); -- 
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652__entry__
      -- CP-element group 4: 	 branch_block_stmt_1642/do_while_stmt_1652/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(4) <= SoftwareRegisterAccessDaemon_CP_2481_elements(3);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	184 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652__exit__
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_back
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	182 
    -- CP-element group 7: 	183 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1642/do_while_stmt_1652/condition_done
      -- CP-element group 7: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_taken/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(7) <= SoftwareRegisterAccessDaemon_CP_2481_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	181 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_body_done
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(8) <= SoftwareRegisterAccessDaemon_CP_2481_elements(181);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	21 
    -- CP-element group 9: 	78 
    -- CP-element group 9: 	59 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/back_edge_to_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(9) <= SoftwareRegisterAccessDaemon_CP_2481_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	42 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	80 
    -- CP-element group 10: 	61 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/first_time_through_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(10) <= SoftwareRegisterAccessDaemon_CP_2481_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	132 
    -- CP-element group 11: 	117 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	108 
    -- CP-element group 11: 	139 
    -- CP-element group 11: 	174 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	73 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	35 
    -- CP-element group 11:  members (12) 
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_root_address_calculated
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	174 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/condition_evaluated
      -- 
    condition_evaluated_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(12), ack => do_while_stmt_1652_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(16) & SoftwareRegisterAccessDaemon_CP_2481_elements(174);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	72 
    -- CP-element group 13: 	53 
    -- CP-element group 13: 	34 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	36 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_sample_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/aggregated_phi_sample_req
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(17) & SoftwareRegisterAccessDaemon_CP_2481_elements(72) & SoftwareRegisterAccessDaemon_CP_2481_elements(53) & SoftwareRegisterAccessDaemon_CP_2481_elements(34) & SoftwareRegisterAccessDaemon_CP_2481_elements(16);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	56 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	181 
    -- CP-element group 14: 	140 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	72 
    -- CP-element group 14: 	53 
    -- CP-element group 14: 	34 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_sample_completed_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(19) & SoftwareRegisterAccessDaemon_CP_2481_elements(37) & SoftwareRegisterAccessDaemon_CP_2481_elements(75) & SoftwareRegisterAccessDaemon_CP_2481_elements(56);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	73 
    -- CP-element group 15: 	54 
    -- CP-element group 15: 	35 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	76 
    -- CP-element group 15: 	57 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_update_start__ps
      -- CP-element group 15: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/aggregated_phi_update_req
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(18) & SoftwareRegisterAccessDaemon_CP_2481_elements(73) & SoftwareRegisterAccessDaemon_CP_2481_elements(54) & SoftwareRegisterAccessDaemon_CP_2481_elements(35);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	77 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/aggregated_phi_update_ack
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(39) & SoftwareRegisterAccessDaemon_CP_2481_elements(77) & SoftwareRegisterAccessDaemon_CP_2481_elements(58);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	123 
    -- CP-element group 18: 	119 
    -- CP-element group 18: 	104 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	100 
    -- CP-element group 18: 	134 
    -- CP-element group 18: 	137 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(123) & SoftwareRegisterAccessDaemon_CP_2481_elements(119) & SoftwareRegisterAccessDaemon_CP_2481_elements(104) & SoftwareRegisterAccessDaemon_CP_2481_elements(97) & SoftwareRegisterAccessDaemon_CP_2481_elements(100) & SoftwareRegisterAccessDaemon_CP_2481_elements(134) & SoftwareRegisterAccessDaemon_CP_2481_elements(137);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: 	132 
    -- CP-element group 20: 	121 
    -- CP-element group 20: 	117 
    -- CP-element group 20: 	95 
    -- CP-element group 20: 	102 
    -- CP-element group 20: 	99 
    -- CP-element group 20: 	136 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(21) <= SoftwareRegisterAccessDaemon_CP_2481_elements(9);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_loopback_sample_req_ps
      -- 
    phi_stmt_1654_loopback_sample_req_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1654_loopback_sample_req_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(22), ack => phi_stmt_1654_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(23) <= SoftwareRegisterAccessDaemon_CP_2481_elements(10);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_entry_sample_req_ps
      -- 
    phi_stmt_1654_entry_sample_req_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1654_entry_sample_req_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(24), ack => phi_stmt_1654_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1654_phi_mux_ack_ps
      -- 
    phi_stmt_1654_phi_mux_ack_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1654_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(28) <= SoftwareRegisterAccessDaemon_CP_2481_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1657_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(27), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_sample_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(32) <= SoftwareRegisterAccessDaemon_CP_2481_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1659_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(31), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	14 
    -- CP-element group 34: 	142 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	13 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(14) & SoftwareRegisterAccessDaemon_CP_2481_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	104 
    -- CP-element group 35: 	97 
    -- CP-element group 35: 	100 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	15 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(104) & SoftwareRegisterAccessDaemon_CP_2481_elements(97) & SoftwareRegisterAccessDaemon_CP_2481_elements(100);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(36) <= SoftwareRegisterAccessDaemon_CP_2481_elements(13);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(38) <= SoftwareRegisterAccessDaemon_CP_2481_elements(15);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: 	95 
    -- CP-element group 39: 	102 
    -- CP-element group 39: 	99 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(40) <= SoftwareRegisterAccessDaemon_CP_2481_elements(9);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_loopback_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_loopback_sample_req
      -- 
    phi_stmt_1660_loopback_sample_req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1660_loopback_sample_req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(41), ack => phi_stmt_1660_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	10 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(42) <= SoftwareRegisterAccessDaemon_CP_2481_elements(10);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_entry_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_entry_sample_req
      -- 
    phi_stmt_1660_entry_sample_req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1660_entry_sample_req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(43), ack => phi_stmt_1660_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_phi_mux_ack_ps
      -- CP-element group 44: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1660_phi_mux_ack
      -- 
    phi_stmt_1660_phi_mux_ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1660_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(47) <= SoftwareRegisterAccessDaemon_CP_2481_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1663_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(46), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_sample_start__ps
      -- 
    req_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(49), ack => check_control_regsiter_1774_1664_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Update/req
      -- CP-element group 50: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_update_start__ps
      -- 
    req_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(50), ack => check_control_regsiter_1774_1664_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_sample_completed__ps
      -- 
    ack_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1774_1664_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_control_regsiter_1664_update_completed__ps
      -- 
    ack_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1774_1664_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	14 
    -- CP-element group 53: 	142 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(14) & SoftwareRegisterAccessDaemon_CP_2481_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	123 
    -- CP-element group 54: 	119 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	15 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(123) & SoftwareRegisterAccessDaemon_CP_2481_elements(119);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(55) <= SoftwareRegisterAccessDaemon_CP_2481_elements(13);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	15 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(57) <= SoftwareRegisterAccessDaemon_CP_2481_elements(15);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	121 
    -- CP-element group 58: 	117 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	9 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(59) <= SoftwareRegisterAccessDaemon_CP_2481_elements(9);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_loopback_sample_req_ps
      -- CP-element group 60: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_loopback_sample_req
      -- 
    phi_stmt_1665_loopback_sample_req_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1665_loopback_sample_req_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(60), ack => phi_stmt_1665_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	10 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(61) <= SoftwareRegisterAccessDaemon_CP_2481_elements(10);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_entry_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_entry_sample_req
      -- 
    phi_stmt_1665_entry_sample_req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1665_entry_sample_req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(62), ack => phi_stmt_1665_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_phi_mux_ack_ps
      -- CP-element group 63: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1665_phi_mux_ack
      -- 
    phi_stmt_1665_phi_mux_ack_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1665_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_sample_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(66) <= SoftwareRegisterAccessDaemon_CP_2481_elements(67);
    -- CP-element group 67:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	66 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1668_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(65), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Sample/req
      -- CP-element group 68: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_sample_start__ps
      -- 
    req_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(68), ack => check_free_q_1783_1669_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Update/req
      -- CP-element group 69: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_update_start_
      -- CP-element group 69: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_update_start__ps
      -- 
    req_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(69), ack => check_free_q_1783_1669_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Sample/ack
      -- CP-element group 70: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_sample_completed__ps
      -- 
    ack_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1783_1669_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Update/ack
      -- CP-element group 71: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_free_q_1669_update_completed__ps
      -- 
    ack_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1783_1669_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	14 
    -- CP-element group 72: 	142 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	13 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(14) & SoftwareRegisterAccessDaemon_CP_2481_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	11 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	134 
    -- CP-element group 73: 	137 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	15 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(134) & SoftwareRegisterAccessDaemon_CP_2481_elements(137);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(74) <= SoftwareRegisterAccessDaemon_CP_2481_elements(13);
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	15 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(76) <= SoftwareRegisterAccessDaemon_CP_2481_elements(15);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	16 
    -- CP-element group 77: 	132 
    -- CP-element group 77: 	136 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(78) <= SoftwareRegisterAccessDaemon_CP_2481_elements(9);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_loopback_sample_req
      -- CP-element group 79: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_loopback_sample_req_ps
      -- 
    phi_stmt_1670_loopback_sample_req_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1670_loopback_sample_req_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(79), ack => phi_stmt_1670_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	10 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(80) <= SoftwareRegisterAccessDaemon_CP_2481_elements(10);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_entry_sample_req_ps
      -- CP-element group 81: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_entry_sample_req
      -- 
    phi_stmt_1670_entry_sample_req_2699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1670_entry_sample_req_2699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(81), ack => phi_stmt_1670_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_phi_mux_ack
      -- CP-element group 82: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/phi_stmt_1670_phi_mux_ack_ps
      -- 
    phi_stmt_1670_phi_mux_ack_2702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1670_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_sample_start__ps
      -- CP-element group 83: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(85) <= SoftwareRegisterAccessDaemon_CP_2481_elements(86);
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	85 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1673_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(84), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_sample_start_
      -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(87), ack => check_num_server_1792_1674_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Update/$entry
      -- 
    req_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(88), ack => check_num_server_1792_1674_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Sample/ack
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1792_1674_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/R_check_num_server_1674_update_completed__ps
      -- 
    ack_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1792_1674_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	11 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	166 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/word_access_start/word_0/rr
      -- CP-element group 91: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/word_access_start/word_0/$entry
      -- 
    rr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(91), ack => array_obj_ref_1679_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(93) & SoftwareRegisterAccessDaemon_CP_2481_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/word_access_complete/$entry
      -- 
    cr_2758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(92), ack => array_obj_ref_1679_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(94);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	175 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/word_access_start/word_0/ra
      -- CP-element group 93: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/word_access_start/$exit
      -- CP-element group 93: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Sample/word_access_start/word_0/$exit
      -- 
    ra_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1679_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	181 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/array_obj_ref_1679_Merge/$entry
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/word_access_complete/word_0/$exit
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/array_obj_ref_1679_Merge/merge_ack
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/word_access_complete/$exit
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/array_obj_ref_1679_Merge/merge_req
      -- CP-element group 94: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_Update/array_obj_ref_1679_Merge/$exit
      -- 
    ca_2759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1679_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	11 
    -- CP-element group 95: 	20 
    -- CP-element group 95: 	39 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	166 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/word_access_start/word_0/rr
      -- CP-element group 95: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/word_access_start/word_0/$entry
      -- CP-element group 95: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/word_access_start/$entry
      -- CP-element group 95: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/$entry
      -- 
    rr_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(95), ack => array_obj_ref_1710_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(39) & SoftwareRegisterAccessDaemon_CP_2481_elements(97) & SoftwareRegisterAccessDaemon_CP_2481_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	100 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/word_access_complete/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_update_start_
      -- CP-element group 96: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/word_access_complete/$entry
      -- CP-element group 96: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/word_access_complete/word_0/cr
      -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(96), ack => array_obj_ref_1710_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(100);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	176 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	35 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Sample/word_access_start/word_0/ra
      -- 
    ra_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1710_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/array_obj_ref_1710_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/array_obj_ref_1710_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/array_obj_ref_1710_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_Update/array_obj_ref_1710_Merge/merge_ack
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1710_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	20 
    -- CP-element group 99: 	39 
    -- CP-element group 99: 	98 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Sample/req
      -- CP-element group 99: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_sample_start_
      -- 
    req_2806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(99), ack => WPIPE_CONTROL_REGISTER_1708_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(39) & SoftwareRegisterAccessDaemon_CP_2481_elements(98) & SoftwareRegisterAccessDaemon_CP_2481_elements(101);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	18 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	35 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Update/req
      -- CP-element group 100: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Sample/ack
      -- CP-element group 100: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_update_start_
      -- 
    ack_2807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1708_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(100)); -- 
    req_2811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(100), ack => WPIPE_CONTROL_REGISTER_1708_inst_req_1); -- 
    -- CP-element group 101:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	181 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	99 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Update/ack
      -- CP-element group 101: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_CONTROL_REGISTER_1708_update_completed_
      -- 
    ack_2812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1708_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(101)); -- 
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: 	39 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Sample/req
      -- 
    req_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(102), ack => W_update_control_register_pipe_1690_delayed_5_0_1712_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(39) & SoftwareRegisterAccessDaemon_CP_2481_elements(104);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	115 
    -- CP-element group 103: 	110 
    -- CP-element group 103: 	112 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_update_start_
      -- CP-element group 103: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Update/req
      -- 
    req_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(103), ack => W_update_control_register_pipe_1690_delayed_5_0_1712_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(115) & SoftwareRegisterAccessDaemon_CP_2481_elements(110) & SoftwareRegisterAccessDaemon_CP_2481_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	18 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	35 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Sample/ack
      -- 
    ack_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_control_register_pipe_1690_delayed_5_0_1712_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(104)); -- 
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	114 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1714_Update/ack
      -- 
    ack_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_control_register_pipe_1690_delayed_5_0_1712_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: 	111 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	112 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	112 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Sample/rr
      -- 
    rr_2868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(106), ack => EQ_u32_u1_1721_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(105) & SoftwareRegisterAccessDaemon_CP_2481_elements(111) & SoftwareRegisterAccessDaemon_CP_2481_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	115 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	113 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Update/cr
      -- 
    cr_2873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(107), ack => EQ_u32_u1_1721_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(115);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	11 
    -- CP-element group 108: 	105 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: 	166 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/word_access_start/$entry
      -- CP-element group 108: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/word_access_start/word_0/rr
      -- 
    rr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(108), ack => array_obj_ref_1718_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(105) & SoftwareRegisterAccessDaemon_CP_2481_elements(110) & SoftwareRegisterAccessDaemon_CP_2481_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	112 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/word_access_complete/$entry
      -- CP-element group 109: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/word_access_complete/word_0/$entry
      -- CP-element group 109: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/word_access_complete/word_0/cr
      -- 
    cr_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(109), ack => array_obj_ref_1718_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	177 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Sample/word_access_start/word_0/ra
      -- 
    ra_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1718_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	106 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/word_access_complete/word_0/ca
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/array_obj_ref_1718_Merge/$entry
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/array_obj_ref_1718_Merge/$exit
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/array_obj_ref_1718_Merge/merge_req
      -- CP-element group 111: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_Update/array_obj_ref_1718_Merge/merge_ack
      -- 
    ca_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1718_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	106 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	103 
    -- CP-element group 112: 	106 
    -- CP-element group 112: 	109 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Sample/ra
      -- 
    ra_2869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_1721_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	107 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/EQ_u32_u1_1721_Update/ca
      -- 
    ca_2874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_1721_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	105 
    -- CP-element group 114: 	113 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Sample/req
      -- 
    req_2882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(114), ack => WPIPE_enable_mac_1716_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(105) & SoftwareRegisterAccessDaemon_CP_2481_elements(113) & SoftwareRegisterAccessDaemon_CP_2481_elements(116);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	103 
    -- CP-element group 115: 	107 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Sample/ack
      -- CP-element group 115: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Update/req
      -- 
    ack_2883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_enable_mac_1716_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(115)); -- 
    req_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(115), ack => WPIPE_enable_mac_1716_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	181 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_enable_mac_1716_Update/ack
      -- 
    ack_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_enable_mac_1716_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	11 
    -- CP-element group 117: 	20 
    -- CP-element group 117: 	58 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	166 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/word_access_start/$entry
      -- CP-element group 117: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/word_access_start/word_0/$entry
      -- CP-element group 117: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/word_access_start/word_0/rr
      -- 
    rr_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(117), ack => array_obj_ref_1726_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(58) & SoftwareRegisterAccessDaemon_CP_2481_elements(119) & SoftwareRegisterAccessDaemon_CP_2481_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	127 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_update_start_
      -- CP-element group 118: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/word_access_complete/$entry
      -- CP-element group 118: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/word_access_complete/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/word_access_complete/word_0/cr
      -- 
    cr_2916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(118), ack => array_obj_ref_1726_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(127);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	178 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	18 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	54 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Sample/word_access_start/word_0/ra
      -- 
    ra_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1726_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	125 
    -- CP-element group 120:  members (9) 
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/array_obj_ref_1726_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/array_obj_ref_1726_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/array_obj_ref_1726_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_Update/array_obj_ref_1726_Merge/merge_ack
      -- 
    ca_2917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1726_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	20 
    -- CP-element group 121: 	58 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Sample/req
      -- 
    req_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(121), ack => W_update_free_q_pipe_1703_delayed_5_0_1728_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(58) & SoftwareRegisterAccessDaemon_CP_2481_elements(123);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	127 
    -- CP-element group 122: 	130 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_update_start_
      -- CP-element group 122: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Update/req
      -- 
    req_2935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(122), ack => W_update_free_q_pipe_1703_delayed_5_0_1728_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(127) & SoftwareRegisterAccessDaemon_CP_2481_elements(130);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	18 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	54 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Sample/ack
      -- 
    ack_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1703_delayed_5_0_1728_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(123)); -- 
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	129 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1730_Update/ack
      -- 
    ack_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1703_delayed_5_0_1728_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	120 
    -- CP-element group 125: 	124 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Sample/rr
      -- 
    rr_2944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(125), ack => type_cast_1734_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(120) & SoftwareRegisterAccessDaemon_CP_2481_elements(124) & SoftwareRegisterAccessDaemon_CP_2481_elements(127);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	130 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Update/cr
      -- 
    cr_2949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(126), ack => type_cast_1734_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(130);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	122 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	118 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Sample/ra
      -- 
    ra_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1734_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/type_cast_1734_Update/ca
      -- 
    ca_2950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1734_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: 	124 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Sample/req
      -- 
    req_2958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(129), ack => WPIPE_FREE_Q_1732_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(128) & SoftwareRegisterAccessDaemon_CP_2481_elements(124) & SoftwareRegisterAccessDaemon_CP_2481_elements(131);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	126 
    -- CP-element group 130: 	122 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_update_start_
      -- CP-element group 130: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Sample/ack
      -- CP-element group 130: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Update/req
      -- 
    ack_2959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1732_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(130)); -- 
    req_2963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(130), ack => WPIPE_FREE_Q_1732_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	181 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_FREE_Q_1732_Update/ack
      -- 
    ack_2964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1732_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	11 
    -- CP-element group 132: 	20 
    -- CP-element group 132: 	77 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	166 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/word_access_start/$entry
      -- CP-element group 132: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/word_access_start/word_0/$entry
      -- CP-element group 132: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/word_access_start/word_0/rr
      -- 
    rr_2981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(132), ack => array_obj_ref_1739_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(77) & SoftwareRegisterAccessDaemon_CP_2481_elements(134) & SoftwareRegisterAccessDaemon_CP_2481_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	137 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/word_access_complete/word_0/cr
      -- 
    cr_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(133), ack => array_obj_ref_1739_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(137);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	179 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	18 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	73 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/word_access_start/$exit
      -- CP-element group 134: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/word_access_start/word_0/$exit
      -- CP-element group 134: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Sample/word_access_start/word_0/ra
      -- 
    ra_2982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1739_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/word_access_complete/$exit
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/word_access_complete/word_0/$exit
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/word_access_complete/word_0/ca
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/array_obj_ref_1739_Merge/$entry
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/array_obj_ref_1739_Merge/$exit
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/array_obj_ref_1739_Merge/merge_req
      -- CP-element group 135: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_Update/array_obj_ref_1739_Merge/merge_ack
      -- 
    ca_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1739_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	20 
    -- CP-element group 136: 	135 
    -- CP-element group 136: 	77 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Sample/req
      -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(136), ack => WPIPE_NUMBER_OF_SERVERS_1737_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(20) & SoftwareRegisterAccessDaemon_CP_2481_elements(135) & SoftwareRegisterAccessDaemon_CP_2481_elements(77) & SoftwareRegisterAccessDaemon_CP_2481_elements(138);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	18 
    -- CP-element group 137: 	133 
    -- CP-element group 137: 	73 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_update_start_
      -- CP-element group 137: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Update/req
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1737_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(137)); -- 
    req_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(137), ack => WPIPE_NUMBER_OF_SERVERS_1737_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	181 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_NUMBER_OF_SERVERS_1737_Update/ack
      -- 
    ack_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1737_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	11 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	142 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Sample/rr
      -- 
    rr_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(139), ack => RPIPE_AFB_NIC_REQUEST_1742_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(11) & SoftwareRegisterAccessDaemon_CP_2481_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	14 
    -- CP-element group 140: 	141 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	161 
    -- CP-element group 140: 	153 
    -- CP-element group 140: 	157 
    -- CP-element group 140: 	145 
    -- CP-element group 140: 	149 
    -- CP-element group 140: 	169 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_update_start_
      -- CP-element group 140: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Update/cr
      -- 
    cr_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(140), ack => RPIPE_AFB_NIC_REQUEST_1742_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(14) & SoftwareRegisterAccessDaemon_CP_2481_elements(141) & SoftwareRegisterAccessDaemon_CP_2481_elements(161) & SoftwareRegisterAccessDaemon_CP_2481_elements(153) & SoftwareRegisterAccessDaemon_CP_2481_elements(157) & SoftwareRegisterAccessDaemon_CP_2481_elements(145) & SoftwareRegisterAccessDaemon_CP_2481_elements(149) & SoftwareRegisterAccessDaemon_CP_2481_elements(169);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	140 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Sample/ra
      -- 
    ra_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1742_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	159 
    -- CP-element group 142: 	151 
    -- CP-element group 142: 	155 
    -- CP-element group 142: 	147 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	167 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: 	72 
    -- CP-element group 142: 	53 
    -- CP-element group 142: 	34 
    -- CP-element group 142:  members (29) 
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/RPIPE_AFB_NIC_REQUEST_1742_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_word_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_root_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_offset_calculated
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_resized_0
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_scaled_0
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_computed_0
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_resize_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_resize_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_resize_0/index_resize_req
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_resize_0/index_resize_ack
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_scale_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_scale_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_scale_0/scale_rename_req
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_index_scale_0/scale_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_final_index_sum_regn/$entry
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_final_index_sum_regn/$exit
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_final_index_sum_regn/req
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_final_index_sum_regn/ack
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_base_plus_offset/$entry
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_base_plus_offset/$exit
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_base_plus_offset/sum_rename_req
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_base_plus_offset/sum_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_word_addrgen/$entry
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_word_addrgen/$exit
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_word_addrgen/root_register_req
      -- CP-element group 142: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_word_addrgen/root_register_ack
      -- 
    ca_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1742_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	166 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/word_access_start/word_0/rr
      -- 
    rr_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(143), ack => array_obj_ref_1795_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(142) & SoftwareRegisterAccessDaemon_CP_2481_elements(166) & SoftwareRegisterAccessDaemon_CP_2481_elements(145);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	165 
    -- CP-element group 144: 	172 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/word_access_complete/$entry
      -- CP-element group 144: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/word_access_complete/word_0/$entry
      -- CP-element group 144: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/word_access_complete/word_0/cr
      -- 
    cr_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(144), ack => array_obj_ref_1795_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(165) & SoftwareRegisterAccessDaemon_CP_2481_elements(172);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	180 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	140 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/word_access_start/$exit
      -- CP-element group 145: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Sample/word_access_start/word_0/ra
      -- 
    ra_3073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1795_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	163 
    -- CP-element group 146: 	171 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/word_access_complete/$exit
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/array_obj_ref_1795_Merge/$entry
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/array_obj_ref_1795_Merge/$exit
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/array_obj_ref_1795_Merge/merge_req
      -- CP-element group 146: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_Update/array_obj_ref_1795_Merge/merge_ack
      -- 
    ca_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1795_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	142 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Sample/req
      -- 
    req_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(147), ack => W_index_1777_delayed_5_0_1797_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(142) & SoftwareRegisterAccessDaemon_CP_2481_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	165 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_update_start_
      -- CP-element group 148: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Update/req
      -- 
    req_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(148), ack => W_index_1777_delayed_5_0_1797_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	140 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Sample/ack
      -- 
    ack_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1777_delayed_5_0_1797_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	163 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1799_Update/ack
      -- 
    ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1777_delayed_5_0_1797_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	142 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Sample/req
      -- 
    req_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(151), ack => W_wdata_1776_delayed_5_0_1800_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(142) & SoftwareRegisterAccessDaemon_CP_2481_elements(153);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	165 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_update_start_
      -- CP-element group 152: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Update/req
      -- 
    req_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(152), ack => W_wdata_1776_delayed_5_0_1800_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: 	140 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Sample/ack
      -- 
    ack_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1776_delayed_5_0_1800_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	163 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1802_Update/ack
      -- 
    ack_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1776_delayed_5_0_1800_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	142 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Sample/req
      -- 
    req_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(155), ack => W_bmask_1774_delayed_5_0_1803_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(142) & SoftwareRegisterAccessDaemon_CP_2481_elements(157);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	165 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_update_start_
      -- CP-element group 156: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Update/req
      -- 
    req_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(156), ack => W_bmask_1774_delayed_5_0_1803_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	140 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Sample/ack
      -- 
    ack_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1774_delayed_5_0_1803_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	163 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1805_Update/ack
      -- 
    ack_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1774_delayed_5_0_1803_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	142 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Sample/req
      -- 
    req_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(159), ack => W_rwbar_1773_delayed_5_0_1806_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(142) & SoftwareRegisterAccessDaemon_CP_2481_elements(161);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	165 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_update_start_
      -- CP-element group 160: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Update/req
      -- 
    req_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(160), ack => W_rwbar_1773_delayed_5_0_1806_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	140 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Sample/ack
      -- 
    ack_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1773_delayed_5_0_1806_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1808_Update/ack
      -- 
    ack_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1773_delayed_5_0_1806_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	175 
    -- CP-element group 163: 	176 
    -- CP-element group 163: 	177 
    -- CP-element group 163: 	178 
    -- CP-element group 163: 	179 
    -- CP-element group 163: 	180 
    -- CP-element group 163: 	158 
    -- CP-element group 163: 	162 
    -- CP-element group 163: 	150 
    -- CP-element group 163: 	154 
    -- CP-element group 163: 	146 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Sample/crr
      -- 
    crr_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(163), ack => call_stmt_1815_call_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(175) & SoftwareRegisterAccessDaemon_CP_2481_elements(176) & SoftwareRegisterAccessDaemon_CP_2481_elements(177) & SoftwareRegisterAccessDaemon_CP_2481_elements(178) & SoftwareRegisterAccessDaemon_CP_2481_elements(179) & SoftwareRegisterAccessDaemon_CP_2481_elements(180) & SoftwareRegisterAccessDaemon_CP_2481_elements(158) & SoftwareRegisterAccessDaemon_CP_2481_elements(162) & SoftwareRegisterAccessDaemon_CP_2481_elements(150) & SoftwareRegisterAccessDaemon_CP_2481_elements(154) & SoftwareRegisterAccessDaemon_CP_2481_elements(146) & SoftwareRegisterAccessDaemon_CP_2481_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_update_start_
      -- CP-element group 164: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Update/ccr
      -- 
    ccr_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(164), ack => call_stmt_1815_call_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	160 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	152 
    -- CP-element group 165: 	156 
    -- CP-element group 165: 	148 
    -- CP-element group 165: 	144 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Sample/cra
      -- 
    cra_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1815_call_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	181 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	91 
    -- CP-element group 166: 	132 
    -- CP-element group 166: 	117 
    -- CP-element group 166: 	95 
    -- CP-element group 166: 	108 
    -- CP-element group 166: 	164 
    -- CP-element group 166: 	143 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/call_stmt_1815_Update/cca
      -- CP-element group 166: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/ring_reenable_memory_space_0
      -- 
    cca_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1815_call_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	142 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Sample/req
      -- 
    req_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(167), ack => W_rwbar_1781_delayed_5_0_1816_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(142) & SoftwareRegisterAccessDaemon_CP_2481_elements(169);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	172 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_update_start_
      -- CP-element group 168: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Update/req
      -- 
    req_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(168), ack => W_rwbar_1781_delayed_5_0_1816_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2481_elements(172);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	140 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Sample/ack
      -- 
    ack_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1781_delayed_5_0_1816_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/assign_stmt_1818_Update/ack
      -- 
    ack_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1781_delayed_5_0_1816_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	146 
    -- CP-element group 171: 	170 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Sample/req
      -- 
    req_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(171), ack => WPIPE_AFB_NIC_RESPONSE_1832_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(146) & SoftwareRegisterAccessDaemon_CP_2481_elements(170) & SoftwareRegisterAccessDaemon_CP_2481_elements(173);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	144 
    -- CP-element group 172: 	168 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_update_start_
      -- CP-element group 172: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Sample/ack
      -- CP-element group 172: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Update/req
      -- 
    ack_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1832_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(172)); -- 
    req_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(172), ack => WPIPE_AFB_NIC_RESPONSE_1832_inst_req_1); -- 
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	181 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/WPIPE_AFB_NIC_RESPONSE_1832_Update/ack
      -- 
    ack_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1832_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(173)); -- 
    -- CP-element group 174:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	11 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	12 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(174) is a control-delay.
    cp_element_174_delay: control_delay_element  generic map(name => " 174_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(11), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(174), clk => clk, reset =>reset);
    -- CP-element group 175:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	93 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	163 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1679_call_stmt_1815_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(175) is a control-delay.
    cp_element_175_delay: control_delay_element  generic map(name => " 175_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(93), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(175), clk => clk, reset =>reset);
    -- CP-element group 176:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	97 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	163 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1710_call_stmt_1815_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(176) is a control-delay.
    cp_element_176_delay: control_delay_element  generic map(name => " 176_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(97), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(176), clk => clk, reset =>reset);
    -- CP-element group 177:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	110 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	163 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1718_call_stmt_1815_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(177) is a control-delay.
    cp_element_177_delay: control_delay_element  generic map(name => " 177_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(110), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(177), clk => clk, reset =>reset);
    -- CP-element group 178:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	119 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	163 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1726_call_stmt_1815_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(178) is a control-delay.
    cp_element_178_delay: control_delay_element  generic map(name => " 178_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(119), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(178), clk => clk, reset =>reset);
    -- CP-element group 179:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	134 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	163 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1739_call_stmt_1815_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(179) is a control-delay.
    cp_element_179_delay: control_delay_element  generic map(name => " 179_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(134), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(179), clk => clk, reset =>reset);
    -- CP-element group 180:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	145 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	163 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/array_obj_ref_1795_call_stmt_1815_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2481_elements(180) is a control-delay.
    cp_element_180_delay: control_delay_element  generic map(name => " 180_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2481_elements(145), ack => SoftwareRegisterAccessDaemon_CP_2481_elements(180), clk => clk, reset =>reset);
    -- CP-element group 181:  join  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	14 
    -- CP-element group 181: 	131 
    -- CP-element group 181: 	116 
    -- CP-element group 181: 	94 
    -- CP-element group 181: 	101 
    -- CP-element group 181: 	166 
    -- CP-element group 181: 	138 
    -- CP-element group 181: 	173 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	8 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1642/do_while_stmt_1652/do_while_stmt_1652_loop_body/$exit
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 31,7 => 31);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2481_elements(14) & SoftwareRegisterAccessDaemon_CP_2481_elements(131) & SoftwareRegisterAccessDaemon_CP_2481_elements(116) & SoftwareRegisterAccessDaemon_CP_2481_elements(94) & SoftwareRegisterAccessDaemon_CP_2481_elements(101) & SoftwareRegisterAccessDaemon_CP_2481_elements(166) & SoftwareRegisterAccessDaemon_CP_2481_elements(138) & SoftwareRegisterAccessDaemon_CP_2481_elements(173);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	7 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_exit/$exit
      -- CP-element group 182: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_exit/ack
      -- 
    ack_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1652_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	7 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_taken/$exit
      -- CP-element group 183: 	 branch_block_stmt_1642/do_while_stmt_1652/loop_taken/ack
      -- 
    ack_3203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1652_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2481_elements(183)); -- 
    -- CP-element group 184:  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	5 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	1 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_1642/do_while_stmt_1652/$exit
      -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(184) <= SoftwareRegisterAccessDaemon_CP_2481_elements(5);
    -- CP-element group 185:  merge  branch  transition  place  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	0 
    -- CP-element group 185: 	2 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	2 
    -- CP-element group 185: 	3 
    -- CP-element group 185:  members (37) 
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_else_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_if_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/merge_stmt_1643__exit__
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646__entry__
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_dead_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/EQ_u1_u1_1649_place
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Sample/req
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Update/cr
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/Update/ca
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/SplitProtocol/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Update/ack
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/branch_req
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Update/req
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/if_stmt_1646_eval_test/EQ_u1_u1_1649/EQ_u1_u1_1649_inputs/RPIPE_MAC_ENABLE_1647/Sample/ack
      -- CP-element group 185: 	 branch_block_stmt_1642/merge_stmt_1643_PhiReqMerge
      -- CP-element group 185: 	 branch_block_stmt_1642/merge_stmt_1643_PhiAck/$entry
      -- CP-element group 185: 	 branch_block_stmt_1642/merge_stmt_1643_PhiAck/$exit
      -- CP-element group 185: 	 branch_block_stmt_1642/merge_stmt_1643_PhiAck/dummy
      -- 
    branch_req_2534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2481_elements(185), ack => if_stmt_1646_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_CP_2481_elements(185) <= OrReduce(SoftwareRegisterAccessDaemon_CP_2481_elements(0) & SoftwareRegisterAccessDaemon_CP_2481_elements(2));
    SoftwareRegisterAccessDaemon_do_while_stmt_1652_terminator_3204: loop_terminator -- 
      generic map (name => " SoftwareRegisterAccessDaemon_do_while_stmt_1652_terminator_3204", max_iterations_in_flight =>31) 
      port map(loop_body_exit => SoftwareRegisterAccessDaemon_CP_2481_elements(8),loop_continue => SoftwareRegisterAccessDaemon_CP_2481_elements(183),loop_terminate => SoftwareRegisterAccessDaemon_CP_2481_elements(182),loop_back => SoftwareRegisterAccessDaemon_CP_2481_elements(6),loop_exit => SoftwareRegisterAccessDaemon_CP_2481_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_1654_phi_seq_2598_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(21);
      SoftwareRegisterAccessDaemon_CP_2481_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(26);
      SoftwareRegisterAccessDaemon_CP_2481_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(28);
      SoftwareRegisterAccessDaemon_CP_2481_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(23);
      SoftwareRegisterAccessDaemon_CP_2481_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(30);
      SoftwareRegisterAccessDaemon_CP_2481_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(32);
      SoftwareRegisterAccessDaemon_CP_2481_elements(24) <= phi_mux_reqs(1);
      phi_stmt_1654_phi_seq_2598 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1654_phi_seq_2598") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2481_elements(13), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(19), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2481_elements(15), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(20), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1660_phi_seq_2642_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(42);
      SoftwareRegisterAccessDaemon_CP_2481_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(45);
      SoftwareRegisterAccessDaemon_CP_2481_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(47);
      SoftwareRegisterAccessDaemon_CP_2481_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(40);
      SoftwareRegisterAccessDaemon_CP_2481_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(51);
      SoftwareRegisterAccessDaemon_CP_2481_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(52);
      SoftwareRegisterAccessDaemon_CP_2481_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1660_phi_seq_2642 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1660_phi_seq_2642") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2481_elements(36), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(37), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2481_elements(38), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(39), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1665_phi_seq_2686_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(61);
      SoftwareRegisterAccessDaemon_CP_2481_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(64);
      SoftwareRegisterAccessDaemon_CP_2481_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(66);
      SoftwareRegisterAccessDaemon_CP_2481_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(59);
      SoftwareRegisterAccessDaemon_CP_2481_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(70);
      SoftwareRegisterAccessDaemon_CP_2481_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(71);
      SoftwareRegisterAccessDaemon_CP_2481_elements(60) <= phi_mux_reqs(1);
      phi_stmt_1665_phi_seq_2686 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1665_phi_seq_2686") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2481_elements(55), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(56), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2481_elements(57), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(58), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1670_phi_seq_2730_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(80);
      SoftwareRegisterAccessDaemon_CP_2481_elements(83)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(83);
      SoftwareRegisterAccessDaemon_CP_2481_elements(84)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(85);
      SoftwareRegisterAccessDaemon_CP_2481_elements(81) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(78);
      SoftwareRegisterAccessDaemon_CP_2481_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(89);
      SoftwareRegisterAccessDaemon_CP_2481_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(90);
      SoftwareRegisterAccessDaemon_CP_2481_elements(79) <= phi_mux_reqs(1);
      phi_stmt_1670_phi_seq_2730 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1670_phi_seq_2730") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2481_elements(74), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(75), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2481_elements(76), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(77), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2481_elements(82), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2560_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(9);
        preds(1)  <= SoftwareRegisterAccessDaemon_CP_2481_elements(10);
        entry_tmerge_2560 : transition_merge -- 
          generic map(name => " entry_tmerge_2560")
          port map (preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2481_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1688_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1696_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1704_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1649_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1772_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1781_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1790_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_1721_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1769_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1778_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1787_wire : std_logic_vector(0 downto 0);
    signal FREE_Q_32_1727 : std_logic_vector(31 downto 0);
    signal INIT_1654 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1685_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1693_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1701_wire : std_logic_vector(0 downto 0);
    signal RPIPE_MAC_ENABLE_1647_wire : std_logic_vector(0 downto 0);
    signal R_index_1794_resized : std_logic_vector(5 downto 0);
    signal R_index_1794_scaled : std_logic_vector(5 downto 0);
    signal addr_1757 : std_logic_vector(35 downto 0);
    signal array_obj_ref_1679_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1679_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1710_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1710_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1710_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1718_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1718_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1718_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1726_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1726_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1739_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1739_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1739_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1795_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1795_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_1795_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1795_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1795_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1795_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1795_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_1753 : std_logic_vector(3 downto 0);
    signal bmask_1774_delayed_5_0_1805 : std_logic_vector(3 downto 0);
    signal check_control_regsiter_1774 : std_logic_vector(0 downto 0);
    signal check_control_regsiter_1774_1664_buffered : std_logic_vector(0 downto 0);
    signal check_free_q_1783 : std_logic_vector(0 downto 0);
    signal check_free_q_1783_1669_buffered : std_logic_vector(0 downto 0);
    signal check_num_server_1792 : std_logic_vector(0 downto 0);
    signal check_num_server_1792_1674_buffered : std_logic_vector(0 downto 0);
    signal control_data_1680 : std_logic_vector(31 downto 0);
    signal control_register_1660 : std_logic_vector(0 downto 0);
    signal free_q_1665 : std_logic_vector(0 downto 0);
    signal index_1765 : std_logic_vector(5 downto 0);
    signal index_1777_delayed_5_0_1799 : std_logic_vector(5 downto 0);
    signal konst_1648_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1768_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1771_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1777_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1780_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1786_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1789_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1836_wire_constant : std_logic_vector(0 downto 0);
    signal num_server_1670 : std_logic_vector(0 downto 0);
    signal rdata_1825 : std_logic_vector(31 downto 0);
    signal req_1743 : std_logic_vector(73 downto 0);
    signal resp_1831 : std_logic_vector(32 downto 0);
    signal rval_1796 : std_logic_vector(31 downto 0);
    signal rwbar_1749 : std_logic_vector(0 downto 0);
    signal rwbar_1773_delayed_5_0_1808 : std_logic_vector(0 downto 0);
    signal rwbar_1781_delayed_5_0_1818 : std_logic_vector(0 downto 0);
    signal type_cast_1657_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1659_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1663_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1668_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1673_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1720_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1734_wire : std_logic_vector(35 downto 0);
    signal type_cast_1823_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1828_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1690 : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1690_delayed_5_0_1714 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1698 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1703_delayed_5_0_1730 : std_logic_vector(0 downto 0);
    signal update_server_num_1706 : std_logic_vector(0 downto 0);
    signal wdata_1761 : std_logic_vector(31 downto 0);
    signal wdata_1776_delayed_5_0_1802 : std_logic_vector(31 downto 0);
    signal wval_1815 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1679_word_address_0 <= "000000";
    array_obj_ref_1710_word_address_0 <= "000000";
    array_obj_ref_1718_word_address_0 <= "000000";
    array_obj_ref_1726_word_address_0 <= "010010";
    array_obj_ref_1739_word_address_0 <= "000001";
    array_obj_ref_1795_offset_scale_factor_0 <= "000001";
    array_obj_ref_1795_resized_base_address <= "000000";
    array_obj_ref_1795_word_offset_0 <= "000000";
    konst_1648_wire_constant <= "0";
    konst_1768_wire_constant <= "000000";
    konst_1771_wire_constant <= "0";
    konst_1777_wire_constant <= "010010";
    konst_1780_wire_constant <= "0";
    konst_1786_wire_constant <= "000001";
    konst_1789_wire_constant <= "0";
    konst_1836_wire_constant <= "1";
    type_cast_1657_wire_constant <= "1";
    type_cast_1659_wire_constant <= "0";
    type_cast_1663_wire_constant <= "0";
    type_cast_1668_wire_constant <= "0";
    type_cast_1673_wire_constant <= "0";
    type_cast_1720_wire_constant <= "00000000000000000000000000000001";
    type_cast_1823_wire_constant <= "00000000000000000000000000000000";
    type_cast_1828_wire_constant <= "0";
    phi_stmt_1654: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1657_wire_constant & type_cast_1659_wire_constant;
      req <= phi_stmt_1654_req_0 & phi_stmt_1654_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1654",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1654_ack_0,
          idata => idata,
          odata => INIT_1654,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1654
    phi_stmt_1660: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1663_wire_constant & check_control_regsiter_1774_1664_buffered;
      req <= phi_stmt_1660_req_0 & phi_stmt_1660_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1660",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1660_ack_0,
          idata => idata,
          odata => control_register_1660,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1660
    phi_stmt_1665: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1668_wire_constant & check_free_q_1783_1669_buffered;
      req <= phi_stmt_1665_req_0 & phi_stmt_1665_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1665",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1665_ack_0,
          idata => idata,
          odata => free_q_1665,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1665
    phi_stmt_1670: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1673_wire_constant & check_num_server_1792_1674_buffered;
      req <= phi_stmt_1670_req_0 & phi_stmt_1670_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1670",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1670_ack_0,
          idata => idata,
          odata => num_server_1670,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1670
    -- flow-through select operator MUX_1824_inst
    rdata_1825 <= rval_1796 when (rwbar_1781_delayed_5_0_1818(0) /=  '0') else type_cast_1823_wire_constant;
    -- flow-through slice operator slice_1748_inst
    rwbar_1749 <= req_1743(72 downto 72);
    -- flow-through slice operator slice_1752_inst
    bmask_1753 <= req_1743(71 downto 68);
    -- flow-through slice operator slice_1756_inst
    addr_1757 <= req_1743(67 downto 32);
    -- flow-through slice operator slice_1760_inst
    wdata_1761 <= req_1743(31 downto 0);
    -- flow-through slice operator slice_1764_inst
    index_1765 <= addr_1757(7 downto 2);
    W_bmask_1774_delayed_5_0_1803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_1774_delayed_5_0_1803_inst_req_0;
      W_bmask_1774_delayed_5_0_1803_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_1774_delayed_5_0_1803_inst_req_1;
      W_bmask_1774_delayed_5_0_1803_inst_ack_1<= rack(0);
      W_bmask_1774_delayed_5_0_1803_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_1774_delayed_5_0_1803_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_1753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_1774_delayed_5_0_1805,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_1777_delayed_5_0_1797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_1777_delayed_5_0_1797_inst_req_0;
      W_index_1777_delayed_5_0_1797_inst_ack_0<= wack(0);
      rreq(0) <= W_index_1777_delayed_5_0_1797_inst_req_1;
      W_index_1777_delayed_5_0_1797_inst_ack_1<= rack(0);
      W_index_1777_delayed_5_0_1797_inst : InterlockBuffer generic map ( -- 
        name => "W_index_1777_delayed_5_0_1797_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_1777_delayed_5_0_1799,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1773_delayed_5_0_1806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1773_delayed_5_0_1806_inst_req_0;
      W_rwbar_1773_delayed_5_0_1806_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1773_delayed_5_0_1806_inst_req_1;
      W_rwbar_1773_delayed_5_0_1806_inst_ack_1<= rack(0);
      W_rwbar_1773_delayed_5_0_1806_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1773_delayed_5_0_1806_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1749,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1773_delayed_5_0_1808,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1781_delayed_5_0_1816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1781_delayed_5_0_1816_inst_req_0;
      W_rwbar_1781_delayed_5_0_1816_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1781_delayed_5_0_1816_inst_req_1;
      W_rwbar_1781_delayed_5_0_1816_inst_ack_1<= rack(0);
      W_rwbar_1781_delayed_5_0_1816_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1781_delayed_5_0_1816_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1749,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1781_delayed_5_0_1818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_control_register_pipe_1690_delayed_5_0_1712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_control_register_pipe_1690_delayed_5_0_1712_inst_req_0;
      W_update_control_register_pipe_1690_delayed_5_0_1712_inst_ack_0<= wack(0);
      rreq(0) <= W_update_control_register_pipe_1690_delayed_5_0_1712_inst_req_1;
      W_update_control_register_pipe_1690_delayed_5_0_1712_inst_ack_1<= rack(0);
      W_update_control_register_pipe_1690_delayed_5_0_1712_inst : InterlockBuffer generic map ( -- 
        name => "W_update_control_register_pipe_1690_delayed_5_0_1712_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_control_register_pipe_1690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_control_register_pipe_1690_delayed_5_0_1714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_free_q_pipe_1703_delayed_5_0_1728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_free_q_pipe_1703_delayed_5_0_1728_inst_req_0;
      W_update_free_q_pipe_1703_delayed_5_0_1728_inst_ack_0<= wack(0);
      rreq(0) <= W_update_free_q_pipe_1703_delayed_5_0_1728_inst_req_1;
      W_update_free_q_pipe_1703_delayed_5_0_1728_inst_ack_1<= rack(0);
      W_update_free_q_pipe_1703_delayed_5_0_1728_inst : InterlockBuffer generic map ( -- 
        name => "W_update_free_q_pipe_1703_delayed_5_0_1728_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_free_q_pipe_1698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_free_q_pipe_1703_delayed_5_0_1730,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_1776_delayed_5_0_1800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_1776_delayed_5_0_1800_inst_req_0;
      W_wdata_1776_delayed_5_0_1800_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_1776_delayed_5_0_1800_inst_req_1;
      W_wdata_1776_delayed_5_0_1800_inst_ack_1<= rack(0);
      W_wdata_1776_delayed_5_0_1800_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_1776_delayed_5_0_1800_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_1761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_1776_delayed_5_0_1802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_control_regsiter_1774_1664_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_control_regsiter_1774_1664_buf_req_0;
      check_control_regsiter_1774_1664_buf_ack_0<= wack(0);
      rreq(0) <= check_control_regsiter_1774_1664_buf_req_1;
      check_control_regsiter_1774_1664_buf_ack_1<= rack(0);
      check_control_regsiter_1774_1664_buf : InterlockBuffer generic map ( -- 
        name => "check_control_regsiter_1774_1664_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_control_regsiter_1774,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_control_regsiter_1774_1664_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_free_q_1783_1669_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_free_q_1783_1669_buf_req_0;
      check_free_q_1783_1669_buf_ack_0<= wack(0);
      rreq(0) <= check_free_q_1783_1669_buf_req_1;
      check_free_q_1783_1669_buf_ack_1<= rack(0);
      check_free_q_1783_1669_buf : InterlockBuffer generic map ( -- 
        name => "check_free_q_1783_1669_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_free_q_1783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_free_q_1783_1669_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_num_server_1792_1674_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_num_server_1792_1674_buf_req_0;
      check_num_server_1792_1674_buf_ack_0<= wack(0);
      rreq(0) <= check_num_server_1792_1674_buf_req_1;
      check_num_server_1792_1674_buf_ack_1<= rack(0);
      check_num_server_1792_1674_buf : InterlockBuffer generic map ( -- 
        name => "check_num_server_1792_1674_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_num_server_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_num_server_1792_1674_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1734_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1734_inst_req_0;
      type_cast_1734_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1734_inst_req_1;
      type_cast_1734_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  update_free_q_pipe_1703_delayed_5_0_1730(0);
      type_cast_1734_inst_gI: SplitGuardInterface generic map(name => "type_cast_1734_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1734_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1734_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => FREE_Q_32_1727,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1734_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1679_gather_scatter
    process(array_obj_ref_1679_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1679_data_0;
      ov(31 downto 0) := iv;
      control_data_1680 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1710_gather_scatter
    process(array_obj_ref_1710_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1710_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1710_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1718_gather_scatter
    process(array_obj_ref_1718_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1718_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1718_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1726_gather_scatter
    process(array_obj_ref_1726_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1726_data_0;
      ov(31 downto 0) := iv;
      FREE_Q_32_1727 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1739_gather_scatter
    process(array_obj_ref_1739_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1739_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1739_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_addr_0
    process(array_obj_ref_1795_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1795_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_1795_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_gather_scatter
    process(array_obj_ref_1795_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1795_data_0;
      ov(31 downto 0) := iv;
      rval_1796 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_index_0_rename
    process(R_index_1794_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1794_resized;
      ov(5 downto 0) := iv;
      R_index_1794_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_index_0_resize
    process(index_1765) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_1765;
      ov(5 downto 0) := iv;
      R_index_1794_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_index_offset
    process(R_index_1794_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1794_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_1795_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1795_root_address_inst
    process(array_obj_ref_1795_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1795_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_1795_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_1652_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1836_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1652_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1652_branch_req_0,
          ack0 => do_while_stmt_1652_branch_ack_0,
          ack1 => do_while_stmt_1652_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1646_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_1649_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1646_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1646_branch_req_0,
          ack0 => if_stmt_1646_branch_ack_0,
          ack1 => if_stmt_1646_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1688_inst
    process(INIT_1654, control_register_1660) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1654, control_register_1660, tmp_var);
      AND_u1_u1_1688_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1696_inst
    process(INIT_1654, free_q_1665) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1654, free_q_1665, tmp_var);
      AND_u1_u1_1696_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1704_inst
    process(INIT_1654, num_server_1670) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1654, num_server_1670, tmp_var);
      AND_u1_u1_1704_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1773_inst
    process(EQ_u6_u1_1769_wire, EQ_u1_u1_1772_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1769_wire, EQ_u1_u1_1772_wire, tmp_var);
      check_control_regsiter_1774 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1782_inst
    process(EQ_u6_u1_1778_wire, EQ_u1_u1_1781_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1778_wire, EQ_u1_u1_1781_wire, tmp_var);
      check_free_q_1783 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1791_inst
    process(EQ_u6_u1_1787_wire, EQ_u1_u1_1790_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1787_wire, EQ_u1_u1_1790_wire, tmp_var);
      check_num_server_1792 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_1830_inst
    process(type_cast_1828_wire_constant, rdata_1825) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1828_wire_constant, rdata_1825, tmp_var);
      resp_1831 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1649_inst
    process(RPIPE_MAC_ENABLE_1647_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(RPIPE_MAC_ENABLE_1647_wire, konst_1648_wire_constant, tmp_var);
      EQ_u1_u1_1649_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1772_inst
    process(rwbar_1749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1749, konst_1771_wire_constant, tmp_var);
      EQ_u1_u1_1772_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1781_inst
    process(rwbar_1749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1749, konst_1780_wire_constant, tmp_var);
      EQ_u1_u1_1781_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1790_inst
    process(rwbar_1749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1749, konst_1789_wire_constant, tmp_var);
      EQ_u1_u1_1790_wire <= tmp_var; --
    end process;
    -- shared split operator group (11) : EQ_u32_u1_1721_inst 
    ApIntEq_group_11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_1718_wire;
      EQ_u32_u1_1721_wire <= data_out(0 downto 0);
      guard_vector(0)  <= update_control_register_pipe_1690_delayed_5_0_1714(0);
      reqL_unguarded(0) <= EQ_u32_u1_1721_inst_req_0;
      EQ_u32_u1_1721_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_1721_inst_req_1;
      EQ_u32_u1_1721_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_11_gI: SplitGuardInterface generic map(name => "ApIntEq_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- binary operator EQ_u6_u1_1769_inst
    process(index_1765) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1765, konst_1768_wire_constant, tmp_var);
      EQ_u6_u1_1769_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1778_inst
    process(index_1765) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1765, konst_1777_wire_constant, tmp_var);
      EQ_u6_u1_1778_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1787_inst
    process(index_1765) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1765, konst_1786_wire_constant, tmp_var);
      EQ_u6_u1_1787_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1685_inst
    process(INIT_1654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1654, tmp_var);
      NOT_u1_u1_1685_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1693_inst
    process(INIT_1654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1654, tmp_var);
      NOT_u1_u1_1693_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1701_inst
    process(INIT_1654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1654, tmp_var);
      NOT_u1_u1_1701_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1689_inst
    process(NOT_u1_u1_1685_wire, AND_u1_u1_1688_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1685_wire, AND_u1_u1_1688_wire, tmp_var);
      update_control_register_pipe_1690 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1697_inst
    process(NOT_u1_u1_1693_wire, AND_u1_u1_1696_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1693_wire, AND_u1_u1_1696_wire, tmp_var);
      update_free_q_pipe_1698 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1705_inst
    process(NOT_u1_u1_1701_wire, AND_u1_u1_1704_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1701_wire, AND_u1_u1_1704_wire, tmp_var);
      update_server_num_1706 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_1739_load_0 array_obj_ref_1726_load_0 array_obj_ref_1795_load_0 array_obj_ref_1718_load_0 array_obj_ref_1710_load_0 array_obj_ref_1679_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 2, 4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 2, 4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => true, 2 => true, 3 => false, 4 => true, 5 => true);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5, 4 => 5, 5 => 5);
      -- 
    begin -- 
      reqL_unguarded(5) <= array_obj_ref_1739_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_1726_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_1795_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1718_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1710_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1679_load_0_req_0;
      array_obj_ref_1739_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_1726_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_1795_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1718_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1710_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1679_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= array_obj_ref_1739_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_1726_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_1795_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1718_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1710_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1679_load_0_req_1;
      array_obj_ref_1739_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_1726_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_1795_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1718_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1710_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1679_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= update_control_register_pipe_1690(0);
      guard_vector(2)  <= update_control_register_pipe_1690_delayed_5_0_1714(0);
      guard_vector(3)  <=  '1';
      guard_vector(4)  <= update_free_q_pipe_1698(0);
      guard_vector(5)  <= update_server_num_1706(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1739_word_address_0 & array_obj_ref_1726_word_address_0 & array_obj_ref_1795_word_address_0 & array_obj_ref_1718_word_address_0 & array_obj_ref_1710_word_address_0 & array_obj_ref_1679_word_address_0;
      array_obj_ref_1739_data_0 <= data_out(191 downto 160);
      array_obj_ref_1726_data_0 <= data_out(159 downto 128);
      array_obj_ref_1795_data_0 <= data_out(127 downto 96);
      array_obj_ref_1718_data_0 <= data_out(95 downto 64);
      array_obj_ref_1710_data_0 <= data_out(63 downto 32);
      array_obj_ref_1679_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_1742_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1742_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_1742_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1742_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_1742_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_1743 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- read from input-signal MAC_ENABLE
    RPIPE_MAC_ENABLE_1647_wire <= MAC_ENABLE;
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_1832_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1832_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_1832_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1832_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_1832_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_1831;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_CONTROL_REGISTER_1708_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1708_inst_req_0;
      WPIPE_CONTROL_REGISTER_1708_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1708_inst_req_1;
      WPIPE_CONTROL_REGISTER_1708_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1690(0);
      data_in <= array_obj_ref_1710_wire;
      CONTROL_REGISTER_write_1_gI: SplitGuardInterface generic map(name => "CONTROL_REGISTER_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      CONTROL_REGISTER_write_1: OutputPortRevised -- 
        generic map ( name => "CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => CONTROL_REGISTER_pipe_write_req(0),
          oack => CONTROL_REGISTER_pipe_write_ack(0),
          odata => CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_FREE_Q_1732_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_FREE_Q_1732_inst_req_0;
      WPIPE_FREE_Q_1732_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_FREE_Q_1732_inst_req_1;
      WPIPE_FREE_Q_1732_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_1703_delayed_5_0_1730(0);
      data_in <= type_cast_1734_wire;
      FREE_Q_write_2_gI: SplitGuardInterface generic map(name => "FREE_Q_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      FREE_Q_write_2: OutputPortRevised -- 
        generic map ( name => "FREE_Q", data_width => 36, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => FREE_Q_pipe_write_req(0),
          oack => FREE_Q_pipe_write_ack(0),
          odata => FREE_Q_pipe_write_data(35 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_NUMBER_OF_SERVERS_1737_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1737_inst_req_0;
      WPIPE_NUMBER_OF_SERVERS_1737_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1737_inst_req_1;
      WPIPE_NUMBER_OF_SERVERS_1737_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_server_num_1706(0);
      data_in <= array_obj_ref_1739_wire;
      NUMBER_OF_SERVERS_write_3_gI: SplitGuardInterface generic map(name => "NUMBER_OF_SERVERS_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NUMBER_OF_SERVERS_write_3: OutputPortRevised -- 
        generic map ( name => "NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_enable_mac_1716_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_enable_mac_1716_inst_req_0;
      WPIPE_enable_mac_1716_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_enable_mac_1716_inst_req_1;
      WPIPE_enable_mac_1716_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1690_delayed_5_0_1714(0);
      data_in <= EQ_u32_u1_1721_wire;
      enable_mac_write_4_gI: SplitGuardInterface generic map(name => "enable_mac_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      enable_mac_write_4: OutputPortRevised -- 
        generic map ( name => "enable_mac", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => enable_mac_pipe_write_req(0),
          oack => enable_mac_pipe_write_ack(0),
          odata => enable_mac_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1815_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1815_call_req_0;
      call_stmt_1815_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1815_call_req_1;
      call_stmt_1815_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_1773_delayed_5_0_1808(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_1774_delayed_5_0_1805 & rval_1796 & wdata_1776_delayed_5_0_1802 & index_1777_delayed_5_0_1799;
      wval_1815 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end SoftwareRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity UpdateRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    bmask : in  std_logic_vector(3 downto 0);
    rval : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    index : in  std_logic_vector(5 downto 0);
    wval : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity UpdateRegister;
architecture UpdateRegister_arch of UpdateRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 74)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal rval_buffer :  std_logic_vector(31 downto 0);
  signal rval_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(5 downto 0);
  signal index_update_enable: Boolean;
  -- output port buffer signals
  signal wval_buffer :  std_logic_vector(31 downto 0);
  signal wval_update_enable: Boolean;
  signal UpdateRegister_CP_34_start: Boolean;
  signal UpdateRegister_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u16_u32_175_inst_req_0 : boolean;
  signal CONCAT_u16_u32_175_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_175_inst_req_1 : boolean;
  signal CONCAT_u16_u32_175_inst_ack_1 : boolean;
  signal array_obj_ref_178_store_0_req_0 : boolean;
  signal array_obj_ref_178_store_0_ack_0 : boolean;
  signal array_obj_ref_178_store_0_req_1 : boolean;
  signal array_obj_ref_178_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "UpdateRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 74) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(3 downto 0) <= bmask;
  bmask_buffer <= in_buffer_data_out(3 downto 0);
  in_buffer_data_in(35 downto 4) <= rval;
  rval_buffer <= in_buffer_data_out(35 downto 4);
  in_buffer_data_in(67 downto 36) <= wdata;
  wdata_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(73 downto 68) <= index;
  index_buffer <= in_buffer_data_out(73 downto 68);
  in_buffer_data_in(tag_length + 73 downto 74) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 73 downto 74);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  UpdateRegister_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "UpdateRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wval_buffer;
  wval <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  UpdateRegister_CP_34: Block -- control-path 
    signal UpdateRegister_CP_34_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    UpdateRegister_CP_34_elements(0) <= UpdateRegister_CP_34_start;
    UpdateRegister_CP_34_symbol <= UpdateRegister_CP_34_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (39) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_sample_start_
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_update_start_
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Sample/rr
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Update/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Update/cr
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_update_start_
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_offset_calculated
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_resized_0
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_computed_0
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/word_access_complete/word_0/cr
      -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_175_inst_req_0); -- 
    cr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_175_inst_req_1); -- 
    cr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => array_obj_ref_178_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_sample_completed_
      -- CP-element group 1: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Sample/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_175_inst_ack_0, ack => UpdateRegister_CP_34_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_update_completed_
      -- CP-element group 2: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Update/$exit
      -- CP-element group 2: 	 assign_stmt_111_to_assign_stmt_180/CONCAT_u16_u32_175_Update/ca
      -- 
    ca_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_175_inst_ack_1, ack => UpdateRegister_CP_34_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_sample_start_
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/array_obj_ref_178_Split/$entry
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/array_obj_ref_178_Split/$exit
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/array_obj_ref_178_Split/split_req
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/array_obj_ref_178_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/word_access_start/word_0/rr
      -- 
    rr_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(3), ack => array_obj_ref_178_store_0_req_0); -- 
    UpdateRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "UpdateRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= UpdateRegister_CP_34_elements(0) & UpdateRegister_CP_34_elements(2);
      gj_UpdateRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => UpdateRegister_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_sample_completed_
      -- CP-element group 4: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Sample/word_access_start/word_0/ra
      -- 
    ra_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_178_store_0_ack_0, ack => UpdateRegister_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_111_to_assign_stmt_180/$exit
      -- CP-element group 5: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_update_completed_
      -- CP-element group 5: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/$exit
      -- CP-element group 5: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_111_to_assign_stmt_180/array_obj_ref_178_Update/word_access_complete/word_0/ca
      -- 
    ca_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_178_store_0_ack_1, ack => UpdateRegister_CP_34_elements(5)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_165_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_174_wire : std_logic_vector(15 downto 0);
    signal MUX_160_wire : std_logic_vector(7 downto 0);
    signal MUX_164_wire : std_logic_vector(7 downto 0);
    signal MUX_169_wire : std_logic_vector(7 downto 0);
    signal MUX_173_wire : std_logic_vector(7 downto 0);
    signal R_index_177_resized : std_logic_vector(5 downto 0);
    signal R_index_177_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_178_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_178_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_178_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_178_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_178_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_178_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_178_word_offset_0 : std_logic_vector(5 downto 0);
    signal b0_111 : std_logic_vector(0 downto 0);
    signal b1_115 : std_logic_vector(0 downto 0);
    signal b2_119 : std_logic_vector(0 downto 0);
    signal b3_123 : std_logic_vector(0 downto 0);
    signal r0_127 : std_logic_vector(7 downto 0);
    signal r1_131 : std_logic_vector(7 downto 0);
    signal r2_135 : std_logic_vector(7 downto 0);
    signal r3_139 : std_logic_vector(7 downto 0);
    signal w0_143 : std_logic_vector(7 downto 0);
    signal w1_147 : std_logic_vector(7 downto 0);
    signal w2_151 : std_logic_vector(7 downto 0);
    signal w3_155 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_178_offset_scale_factor_0 <= "000001";
    array_obj_ref_178_resized_base_address <= "000000";
    array_obj_ref_178_word_offset_0 <= "000000";
    -- flow-through select operator MUX_160_inst
    MUX_160_wire <= w0_143 when (b0_111(0) /=  '0') else r0_127;
    -- flow-through select operator MUX_164_inst
    MUX_164_wire <= w1_147 when (b1_115(0) /=  '0') else r1_131;
    -- flow-through select operator MUX_169_inst
    MUX_169_wire <= w2_151 when (b2_119(0) /=  '0') else r2_135;
    -- flow-through select operator MUX_173_inst
    MUX_173_wire <= w3_155 when (b3_123(0) /=  '0') else r3_139;
    -- flow-through slice operator slice_110_inst
    b0_111 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_114_inst
    b1_115 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_118_inst
    b2_119 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_122_inst
    b3_123 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_126_inst
    r0_127 <= rval_buffer(31 downto 24);
    -- flow-through slice operator slice_130_inst
    r1_131 <= rval_buffer(23 downto 16);
    -- flow-through slice operator slice_134_inst
    r2_135 <= rval_buffer(15 downto 8);
    -- flow-through slice operator slice_138_inst
    r3_139 <= rval_buffer(7 downto 0);
    -- flow-through slice operator slice_142_inst
    w0_143 <= wdata_buffer(31 downto 24);
    -- flow-through slice operator slice_146_inst
    w1_147 <= wdata_buffer(23 downto 16);
    -- flow-through slice operator slice_150_inst
    w2_151 <= wdata_buffer(15 downto 8);
    -- flow-through slice operator slice_154_inst
    w3_155 <= wdata_buffer(7 downto 0);
    -- equivalence array_obj_ref_178_addr_0
    process(array_obj_ref_178_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_178_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_178_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_178_gather_scatter
    process(wval_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_178_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_178_index_0_rename
    process(R_index_177_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_177_resized;
      ov(5 downto 0) := iv;
      R_index_177_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_178_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(5 downto 0) := iv;
      R_index_177_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_178_index_offset
    process(R_index_177_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_177_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_178_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_178_root_address_inst
    process(array_obj_ref_178_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_178_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_178_root_address <= ov(5 downto 0);
      --
    end process;
    -- shared split operator group (0) : CONCAT_u16_u32_175_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_165_wire & CONCAT_u8_u16_174_wire;
      wval_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_175_inst_req_0;
      CONCAT_u16_u32_175_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_175_inst_req_1;
      CONCAT_u16_u32_175_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u8_u16_165_inst
    process(MUX_160_wire, MUX_164_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_160_wire, MUX_164_wire, tmp_var);
      CONCAT_u8_u16_165_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_174_inst
    process(MUX_169_wire, MUX_173_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_169_wire, MUX_173_wire, tmp_var);
      CONCAT_u8_u16_174_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_178_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_178_store_0_req_0;
      array_obj_ref_178_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_178_store_0_req_1;
      array_obj_ref_178_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_178_word_address_0;
      data_in <= array_obj_ref_178_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(5 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end UpdateRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity accessMemory is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemory;
architecture accessMemory_arch of accessMemory is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 110)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal bmask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemory_CP_513_start: Boolean;
  signal accessMemory_CP_513_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_298_branch_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_ack_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_ack_1 : boolean;
  signal do_while_stmt_298_branch_ack_0 : boolean;
  signal do_while_stmt_298_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemory_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 110) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= bmask;
  bmask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(45 downto 10) <= addr;
  addr_buffer <= in_buffer_data_out(45 downto 10);
  in_buffer_data_in(109 downto 46) <= wdata;
  wdata_buffer <= in_buffer_data_out(109 downto 46);
  in_buffer_data_in(tag_length + 109 downto 110) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 109 downto 110);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemory_CP_513_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemory_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_513_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemory_CP_513_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_513_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemory_CP_513: Block -- control-path 
    signal accessMemory_CP_513_elements: BooleanArray(20 downto 0);
    -- 
  begin -- 
    accessMemory_CP_513_elements(0) <= accessMemory_CP_513_start;
    accessMemory_CP_513_symbol <= accessMemory_CP_513_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_297/$entry
      -- CP-element group 0: 	 branch_block_stmt_297/branch_block_stmt_297__entry__
      -- CP-element group 0: 	 branch_block_stmt_297/do_while_stmt_298__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_297/$exit
      -- CP-element group 1: 	 branch_block_stmt_297/branch_block_stmt_297__exit__
      -- CP-element group 1: 	 branch_block_stmt_297/do_while_stmt_298__exit__
      -- 
    accessMemory_CP_513_elements(1) <= accessMemory_CP_513_elements(20);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_297/do_while_stmt_298/$entry
      -- CP-element group 2: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298__entry__
      -- 
    accessMemory_CP_513_elements(2) <= accessMemory_CP_513_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	20 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298__exit__
      -- 
    -- Element group accessMemory_CP_513_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_297/do_while_stmt_298/loop_back
      -- 
    -- Element group accessMemory_CP_513_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	18 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_297/do_while_stmt_298/condition_done
      -- CP-element group 5: 	 branch_block_stmt_297/do_while_stmt_298/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_297/do_while_stmt_298/loop_taken/$entry
      -- 
    accessMemory_CP_513_elements(5) <= accessMemory_CP_513_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	13 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_297/do_while_stmt_298/loop_body_done
      -- 
    accessMemory_CP_513_elements(6) <= accessMemory_CP_513_elements(13);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/back_edge_to_loop_body
      -- 
    accessMemory_CP_513_elements(7) <= accessMemory_CP_513_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/first_time_through_loop_body
      -- 
    accessMemory_CP_513_elements(8) <= accessMemory_CP_513_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	17 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/loop_body_start
      -- 
    -- Element group accessMemory_CP_513_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	17 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/condition_evaluated
      -- 
    condition_evaluated_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_513_elements(10), ack => do_while_stmt_298_branch_req_0); -- 
    accessMemory_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_513_elements(16) & accessMemory_CP_513_elements(17);
      gj_accessMemory_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_513_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Sample/req
      -- 
    req_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_513_elements(11), ack => WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_req_0); -- 
    accessMemory_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_513_elements(9) & accessMemory_CP_513_elements(13);
      gj_accessMemory_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_513_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_update_start_
      -- CP-element group 12: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Sample/ack
      -- CP-element group 12: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Update/req
      -- 
    ack_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_ack_0, ack => accessMemory_CP_513_elements(12)); -- 
    req_551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_513_elements(12), ack => WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_req_1); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	6 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/$exit
      -- CP-element group 13: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_311_Update/ack
      -- 
    ack_552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_ack_1, ack => accessMemory_CP_513_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Sample/rr
      -- 
    rr_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_513_elements(14), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_req_0); -- 
    accessMemory_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_513_elements(9) & accessMemory_CP_513_elements(16);
      gj_accessMemory_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_513_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_update_start_
      -- CP-element group 15: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Update/cr
      -- 
    ra_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_ack_0, ack => accessMemory_CP_513_elements(15)); -- 
    cr_565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_513_elements(15), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_req_1); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_315_Update/ca
      -- 
    ca_566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_ack_1, ack => accessMemory_CP_513_elements(16)); -- 
    -- CP-element group 17:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	10 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_297/do_while_stmt_298/do_while_stmt_298_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group accessMemory_CP_513_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => accessMemory_CP_513_elements(9), ack => accessMemory_CP_513_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	5 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_297/do_while_stmt_298/loop_exit/$exit
      -- CP-element group 18: 	 branch_block_stmt_297/do_while_stmt_298/loop_exit/ack
      -- 
    ack_571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_298_branch_ack_0, ack => accessMemory_CP_513_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_297/do_while_stmt_298/loop_taken/$exit
      -- CP-element group 19: 	 branch_block_stmt_297/do_while_stmt_298/loop_taken/ack
      -- 
    ack_575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_298_branch_ack_1, ack => accessMemory_CP_513_elements(19)); -- 
    -- CP-element group 20:  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	3 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	1 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_297/do_while_stmt_298/$exit
      -- 
    accessMemory_CP_513_elements(20) <= accessMemory_CP_513_elements(3);
    accessMemory_do_while_stmt_298_terminator_576: loop_terminator -- 
      generic map (name => " accessMemory_do_while_stmt_298_terminator_576", max_iterations_in_flight =>15) 
      port map(loop_body_exit => accessMemory_CP_513_elements(6),loop_continue => accessMemory_CP_513_elements(19),loop_terminate => accessMemory_CP_513_elements(18),loop_back => accessMemory_CP_513_elements(4),loop_exit => accessMemory_CP_513_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_538_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= accessMemory_CP_513_elements(7);
        preds(1)  <= accessMemory_CP_513_elements(8);
        entry_tmerge_538 : transition_merge -- 
          generic map(name => " entry_tmerge_538")
          port map (preds => preds, symbol_out => accessMemory_CP_513_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_303_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_305_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_308_wire : std_logic_vector(99 downto 0);
    signal EQ_u1_u1_334_wire : std_logic_vector(0 downto 0);
    signal err_320 : std_logic_vector(0 downto 0);
    signal konst_333_wire_constant : std_logic_vector(0 downto 0);
    signal request_310 : std_logic_vector(109 downto 0);
    signal response_316 : std_logic_vector(64 downto 0);
    -- 
  begin -- 
    konst_333_wire_constant <= "1";
    -- flow-through slice operator slice_319_inst
    err_320 <= response_316(64 downto 64);
    -- flow-through slice operator slice_323_inst
    rdata_buffer <= response_316(63 downto 0);
    do_while_stmt_298_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_334_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_298_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_298_branch_req_0,
          ack0 => do_while_stmt_298_branch_ack_0,
          ack1 => do_while_stmt_298_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u10_u110_309_inst
    process(CONCAT_u2_u10_305_wire, CONCAT_u36_u100_308_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_305_wire, CONCAT_u36_u100_308_wire, tmp_var);
      request_310 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_303_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_303_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_305_inst
    process(CONCAT_u1_u2_303_wire, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_303_wire, bmask_buffer, tmp_var);
      CONCAT_u2_u10_305_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_308_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_308_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_334_inst
    process(err_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(err_320, konst_333_wire_constant, tmp_var);
      EQ_u1_u1_334_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_315_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_316 <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_TO_MEMORY_REQUEST_311_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_311_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_310;
      NIC_TO_MEMORY_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemory_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity acquireLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireLock;
architecture acquireLock_arch of acquireLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireLock_CP_577_start: Boolean;
  signal acquireLock_CP_577_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_497_branch_req_0 : boolean;
  signal call_stmt_514_call_ack_0 : boolean;
  signal call_stmt_587_call_ack_1 : boolean;
  signal call_stmt_587_call_req_1 : boolean;
  signal call_stmt_587_call_ack_0 : boolean;
  signal call_stmt_514_call_req_0 : boolean;
  signal call_stmt_359_call_req_0 : boolean;
  signal call_stmt_587_call_req_0 : boolean;
  signal call_stmt_359_call_ack_0 : boolean;
  signal call_stmt_359_call_ack_1 : boolean;
  signal call_stmt_383_call_ack_1 : boolean;
  signal call_stmt_383_call_req_1 : boolean;
  signal call_stmt_383_call_ack_0 : boolean;
  signal call_stmt_359_call_req_1 : boolean;
  signal call_stmt_383_call_req_0 : boolean;
  signal if_stmt_497_branch_ack_0 : boolean;
  signal if_stmt_497_branch_ack_1 : boolean;
  signal call_stmt_514_call_ack_1 : boolean;
  signal call_stmt_514_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireLock_CP_577_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_577_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireLock_CP_577_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_577_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireLock_CP_577: Block -- control-path 
    signal acquireLock_CP_577_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    acquireLock_CP_577_elements(0) <= acquireLock_CP_577_start;
    acquireLock_CP_577_symbol <= acquireLock_CP_577_elements(10);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_340/merge_stmt_347__entry__
      -- CP-element group 0: 	 branch_block_stmt_340/merge_stmt_347_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_340/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_340/assign_stmt_346__exit__
      -- CP-element group 0: 	 branch_block_stmt_340/assign_stmt_346__entry__
      -- CP-element group 0: 	 branch_block_stmt_340/merge_stmt_347__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_340/merge_stmt_347__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_340/branch_block_stmt_340__entry__
      -- CP-element group 0: 	 branch_block_stmt_340/assign_stmt_346/$exit
      -- CP-element group 0: 	 branch_block_stmt_340/assign_stmt_346/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	11 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_sample_completed_
      -- 
    cra_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_359_call_ack_0, ack => acquireLock_CP_577_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_sample_start_
      -- 
    cca_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_359_call_ack_1, ack => acquireLock_CP_577_elements(2)); -- 
    crr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(2), ack => call_stmt_383_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_sample_completed_
      -- 
    cra_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_383_call_ack_0, ack => acquireLock_CP_577_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	11 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497__entry__
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/EQ_u8_u1_502_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/EQ_u8_u1_502_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496__exit__
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/EQ_u8_u1_502/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_340/EQ_u8_u1_502_place
      -- CP-element group 4: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/$exit
      -- CP-element group 4: 	 branch_block_stmt_340/if_stmt_497_else_link/$entry
      -- 
    cca_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_383_call_ack_1, ack => acquireLock_CP_577_elements(4)); -- 
    branch_req_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(4), ack => if_stmt_497_branch_req_0); -- 
    -- CP-element group 5:  fork  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (10) 
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Sample/crr
      -- CP-element group 5: 	 branch_block_stmt_340/if_stmt_497_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_update_start_
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/$entry
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514__entry__
      -- CP-element group 5: 	 branch_block_stmt_340/if_stmt_497_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Update/ccr
      -- 
    if_choice_transition_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_497_branch_ack_1, ack => acquireLock_CP_577_elements(5)); -- 
    crr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(5), ack => call_stmt_514_call_req_0); -- 
    ccr_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(5), ack => call_stmt_514_call_req_1); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: 	10 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587__entry__
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Update/ccr
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_update_start_
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/$entry
      -- CP-element group 6: 	 branch_block_stmt_340/if_stmt_497__exit__
      -- CP-element group 6: 	 branch_block_stmt_340/if_stmt_497_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_340/if_stmt_497_else_link/$exit
      -- 
    else_choice_transition_664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_497_branch_ack_0, ack => acquireLock_CP_577_elements(6)); -- 
    ccr_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(6), ack => call_stmt_587_call_req_1); -- 
    crr_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(6), ack => call_stmt_587_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Sample/cra
      -- CP-element group 7: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_sample_completed_
      -- 
    cra_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_514_call_ack_0, ack => acquireLock_CP_577_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (8) 
      -- CP-element group 8: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_340/call_stmt_514/$exit
      -- CP-element group 8: 	 branch_block_stmt_340/loopback
      -- CP-element group 8: 	 branch_block_stmt_340/call_stmt_514__exit__
      -- CP-element group 8: 	 branch_block_stmt_340/loopback_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_340/loopback_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_340/call_stmt_514/call_stmt_514_Update/cca
      -- 
    cca_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_514_call_ack_1, ack => acquireLock_CP_577_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Sample/cra
      -- CP-element group 9: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_sample_completed_
      -- 
    cra_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_587_call_ack_0, ack => acquireLock_CP_577_elements(9)); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	6 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Update/cca
      -- CP-element group 10: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/call_stmt_587_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587/$exit
      -- CP-element group 10: 	 assign_stmt_592/$exit
      -- CP-element group 10: 	 assign_stmt_592/$entry
      -- CP-element group 10: 	 branch_block_stmt_340/$exit
      -- CP-element group 10: 	 $exit
      -- CP-element group 10: 	 branch_block_stmt_340/branch_block_stmt_340__exit__
      -- CP-element group 10: 	 branch_block_stmt_340/assign_stmt_573_to_call_stmt_587__exit__
      -- 
    cca_701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_587_call_ack_1, ack => acquireLock_CP_577_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: 	2 
    -- CP-element group 11: 	4 
    -- CP-element group 11:  members (16) 
      -- CP-element group 11: 	 branch_block_stmt_340/merge_stmt_347_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_340/merge_stmt_347_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Sample/crr
      -- CP-element group 11: 	 branch_block_stmt_340/merge_stmt_347_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_update_start_
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496__entry__
      -- CP-element group 11: 	 branch_block_stmt_340/merge_stmt_347__exit__
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Update/ccr
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_Update/ccr
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_359_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_340/merge_stmt_347_PhiAck/dummy
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/$entry
      -- CP-element group 11: 	 branch_block_stmt_340/call_stmt_359_to_assign_stmt_496/call_stmt_383_update_start_
      -- 
    crr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(11), ack => call_stmt_359_call_req_0); -- 
    ccr_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(11), ack => call_stmt_383_call_req_1); -- 
    ccr_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_577_elements(11), ack => call_stmt_359_call_req_1); -- 
    acquireLock_CP_577_elements(11) <= OrReduce(acquireLock_CP_577_elements(0) & acquireLock_CP_577_elements(8));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_530_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_543_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_557_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_570_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_544_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_571_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u4_u36_379_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u4_u36_582_wire : std_logic_vector(35 downto 0);
    signal EQ_u8_u1_502_wire : std_logic_vector(0 downto 0);
    signal MUX_460_wire : std_logic_vector(7 downto 0);
    signal MUX_464_wire : std_logic_vector(7 downto 0);
    signal MUX_469_wire : std_logic_vector(7 downto 0);
    signal MUX_473_wire : std_logic_vector(7 downto 0);
    signal MUX_479_wire : std_logic_vector(7 downto 0);
    signal MUX_483_wire : std_logic_vector(7 downto 0);
    signal MUX_488_wire : std_logic_vector(7 downto 0);
    signal MUX_492_wire : std_logic_vector(7 downto 0);
    signal MUX_523_wire : std_logic_vector(0 downto 0);
    signal MUX_529_wire : std_logic_vector(0 downto 0);
    signal MUX_536_wire : std_logic_vector(0 downto 0);
    signal MUX_542_wire : std_logic_vector(0 downto 0);
    signal MUX_550_wire : std_logic_vector(0 downto 0);
    signal MUX_556_wire : std_logic_vector(0 downto 0);
    signal MUX_563_wire : std_logic_vector(0 downto 0);
    signal MUX_569_wire : std_logic_vector(0 downto 0);
    signal NOT_u64_u64_585_wire_constant : std_logic_vector(63 downto 0);
    signal NOT_u8_u8_354_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_375_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_501_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_509_wire_constant : std_logic_vector(7 downto 0);
    signal OR_u8_u8_465_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_474_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_475_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_484_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_493_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_494_wire : std_logic_vector(7 downto 0);
    signal err_514 : std_logic_vector(63 downto 0);
    signal ignore_587 : std_logic_vector(63 downto 0);
    signal konst_418_wire_constant : std_logic_vector(2 downto 0);
    signal konst_423_wire_constant : std_logic_vector(2 downto 0);
    signal konst_428_wire_constant : std_logic_vector(2 downto 0);
    signal konst_433_wire_constant : std_logic_vector(2 downto 0);
    signal konst_438_wire_constant : std_logic_vector(2 downto 0);
    signal konst_443_wire_constant : std_logic_vector(2 downto 0);
    signal konst_448_wire_constant : std_logic_vector(2 downto 0);
    signal konst_453_wire_constant : std_logic_vector(2 downto 0);
    signal konst_459_wire_constant : std_logic_vector(7 downto 0);
    signal konst_463_wire_constant : std_logic_vector(7 downto 0);
    signal konst_468_wire_constant : std_logic_vector(7 downto 0);
    signal konst_472_wire_constant : std_logic_vector(7 downto 0);
    signal konst_478_wire_constant : std_logic_vector(7 downto 0);
    signal konst_482_wire_constant : std_logic_vector(7 downto 0);
    signal konst_487_wire_constant : std_logic_vector(7 downto 0);
    signal konst_491_wire_constant : std_logic_vector(7 downto 0);
    signal l0_387 : std_logic_vector(7 downto 0);
    signal l1_391 : std_logic_vector(7 downto 0);
    signal l2_395 : std_logic_vector(7 downto 0);
    signal l3_399 : std_logic_vector(7 downto 0);
    signal l4_403 : std_logic_vector(7 downto 0);
    signal l5_407 : std_logic_vector(7 downto 0);
    signal l6_411 : std_logic_vector(7 downto 0);
    signal l7_415 : std_logic_vector(7 downto 0);
    signal lock_addr_32_363 : std_logic_vector(31 downto 0);
    signal lock_address_pointer_346 : std_logic_vector(35 downto 0);
    signal lock_val_496 : std_logic_vector(7 downto 0);
    signal lock_values_383 : std_logic_vector(63 downto 0);
    signal msg_size_plus_lock_359 : std_logic_vector(63 downto 0);
    signal new_bmask_573 : std_logic_vector(7 downto 0);
    signal s0_420 : std_logic_vector(0 downto 0);
    signal s1_425 : std_logic_vector(0 downto 0);
    signal s2_430 : std_logic_vector(0 downto 0);
    signal s3_435 : std_logic_vector(0 downto 0);
    signal s4_440 : std_logic_vector(0 downto 0);
    signal s5_445 : std_logic_vector(0 downto 0);
    signal s6_450 : std_logic_vector(0 downto 0);
    signal s7_455 : std_logic_vector(0 downto 0);
    signal sel_368 : std_logic_vector(2 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_349_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_351_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_357_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_370_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_372_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_377_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_381_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_504_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_506_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_522_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_526_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_528_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_533_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_535_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_539_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_541_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_549_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_555_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_560_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_562_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_568_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_575_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_577_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_580_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    NOT_u64_u64_585_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    NOT_u8_u8_354_wire_constant <= "11111111";
    NOT_u8_u8_375_wire_constant <= "11111111";
    NOT_u8_u8_501_wire_constant <= "11111111";
    NOT_u8_u8_509_wire_constant <= "11111111";
    konst_418_wire_constant <= "000";
    konst_423_wire_constant <= "001";
    konst_428_wire_constant <= "010";
    konst_433_wire_constant <= "011";
    konst_438_wire_constant <= "100";
    konst_443_wire_constant <= "101";
    konst_448_wire_constant <= "110";
    konst_453_wire_constant <= "111";
    konst_459_wire_constant <= "00000000";
    konst_463_wire_constant <= "00000000";
    konst_468_wire_constant <= "00000000";
    konst_472_wire_constant <= "00000000";
    konst_478_wire_constant <= "00000000";
    konst_482_wire_constant <= "00000000";
    konst_487_wire_constant <= "00000000";
    konst_491_wire_constant <= "00000000";
    type_cast_344_wire_constant <= "000000000000000000000000000000010000";
    type_cast_349_wire_constant <= "1";
    type_cast_351_wire_constant <= "1";
    type_cast_357_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_370_wire_constant <= "1";
    type_cast_372_wire_constant <= "1";
    type_cast_377_wire_constant <= "0000";
    type_cast_381_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_504_wire_constant <= "0";
    type_cast_506_wire_constant <= "1";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_520_wire_constant <= "1";
    type_cast_522_wire_constant <= "0";
    type_cast_526_wire_constant <= "1";
    type_cast_528_wire_constant <= "0";
    type_cast_533_wire_constant <= "1";
    type_cast_535_wire_constant <= "0";
    type_cast_539_wire_constant <= "1";
    type_cast_541_wire_constant <= "0";
    type_cast_547_wire_constant <= "1";
    type_cast_549_wire_constant <= "0";
    type_cast_553_wire_constant <= "1";
    type_cast_555_wire_constant <= "0";
    type_cast_560_wire_constant <= "1";
    type_cast_562_wire_constant <= "0";
    type_cast_566_wire_constant <= "1";
    type_cast_568_wire_constant <= "0";
    type_cast_575_wire_constant <= "0";
    type_cast_577_wire_constant <= "0";
    type_cast_580_wire_constant <= "0000";
    -- flow-through select operator MUX_460_inst
    MUX_460_wire <= l0_387 when (s0_420(0) /=  '0') else konst_459_wire_constant;
    -- flow-through select operator MUX_464_inst
    MUX_464_wire <= l1_391 when (s1_425(0) /=  '0') else konst_463_wire_constant;
    -- flow-through select operator MUX_469_inst
    MUX_469_wire <= l2_395 when (s2_430(0) /=  '0') else konst_468_wire_constant;
    -- flow-through select operator MUX_473_inst
    MUX_473_wire <= l3_399 when (s3_435(0) /=  '0') else konst_472_wire_constant;
    -- flow-through select operator MUX_479_inst
    MUX_479_wire <= l4_403 when (s4_440(0) /=  '0') else konst_478_wire_constant;
    -- flow-through select operator MUX_483_inst
    MUX_483_wire <= l5_407 when (s5_445(0) /=  '0') else konst_482_wire_constant;
    -- flow-through select operator MUX_488_inst
    MUX_488_wire <= l6_411 when (s6_450(0) /=  '0') else konst_487_wire_constant;
    -- flow-through select operator MUX_492_inst
    MUX_492_wire <= l7_415 when (s7_455(0) /=  '0') else konst_491_wire_constant;
    -- flow-through select operator MUX_523_inst
    MUX_523_wire <= type_cast_520_wire_constant when (s0_420(0) /=  '0') else type_cast_522_wire_constant;
    -- flow-through select operator MUX_529_inst
    MUX_529_wire <= type_cast_526_wire_constant when (s1_425(0) /=  '0') else type_cast_528_wire_constant;
    -- flow-through select operator MUX_536_inst
    MUX_536_wire <= type_cast_533_wire_constant when (s2_430(0) /=  '0') else type_cast_535_wire_constant;
    -- flow-through select operator MUX_542_inst
    MUX_542_wire <= type_cast_539_wire_constant when (s3_435(0) /=  '0') else type_cast_541_wire_constant;
    -- flow-through select operator MUX_550_inst
    MUX_550_wire <= type_cast_547_wire_constant when (s4_440(0) /=  '0') else type_cast_549_wire_constant;
    -- flow-through select operator MUX_556_inst
    MUX_556_wire <= type_cast_553_wire_constant when (s5_445(0) /=  '0') else type_cast_555_wire_constant;
    -- flow-through select operator MUX_563_inst
    MUX_563_wire <= type_cast_560_wire_constant when (s6_450(0) /=  '0') else type_cast_562_wire_constant;
    -- flow-through select operator MUX_569_inst
    MUX_569_wire <= type_cast_566_wire_constant when (s7_455(0) /=  '0') else type_cast_568_wire_constant;
    -- flow-through slice operator slice_362_inst
    lock_addr_32_363 <= msg_size_plus_lock_359(31 downto 0);
    -- flow-through slice operator slice_367_inst
    sel_368 <= lock_addr_32_363(2 downto 0);
    -- flow-through slice operator slice_386_inst
    l0_387 <= lock_values_383(63 downto 56);
    -- flow-through slice operator slice_390_inst
    l1_391 <= lock_values_383(55 downto 48);
    -- flow-through slice operator slice_394_inst
    l2_395 <= lock_values_383(47 downto 40);
    -- flow-through slice operator slice_398_inst
    l3_399 <= lock_values_383(39 downto 32);
    -- flow-through slice operator slice_402_inst
    l4_403 <= lock_values_383(31 downto 24);
    -- flow-through slice operator slice_406_inst
    l5_407 <= lock_values_383(23 downto 16);
    -- flow-through slice operator slice_410_inst
    l6_411 <= lock_values_383(15 downto 8);
    -- flow-through slice operator slice_414_inst
    l7_415 <= lock_values_383(7 downto 0);
    if_stmt_497_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u8_u1_502_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_497_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_497_branch_req_0,
          ack0 => if_stmt_497_branch_ack_0,
          ack1 => if_stmt_497_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u36_u36_345_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_344_wire_constant, tmp_var);
      lock_address_pointer_346 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_530_inst
    process(MUX_523_wire, MUX_529_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_523_wire, MUX_529_wire, tmp_var);
      CONCAT_u1_u2_530_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_543_inst
    process(MUX_536_wire, MUX_542_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_536_wire, MUX_542_wire, tmp_var);
      CONCAT_u1_u2_543_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_557_inst
    process(MUX_550_wire, MUX_556_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_550_wire, MUX_556_wire, tmp_var);
      CONCAT_u1_u2_557_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_570_inst
    process(MUX_563_wire, MUX_569_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_563_wire, MUX_569_wire, tmp_var);
      CONCAT_u1_u2_570_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_544_inst
    process(CONCAT_u1_u2_530_wire, CONCAT_u1_u2_543_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_530_wire, CONCAT_u1_u2_543_wire, tmp_var);
      CONCAT_u2_u4_544_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_571_inst
    process(CONCAT_u1_u2_557_wire, CONCAT_u1_u2_570_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_557_wire, CONCAT_u1_u2_570_wire, tmp_var);
      CONCAT_u2_u4_571_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_379_inst
    process(type_cast_377_wire_constant, lock_addr_32_363) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_377_wire_constant, lock_addr_32_363, tmp_var);
      CONCAT_u4_u36_379_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_582_inst
    process(type_cast_580_wire_constant, lock_addr_32_363) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_580_wire_constant, lock_addr_32_363, tmp_var);
      CONCAT_u4_u36_582_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_572_inst
    process(CONCAT_u2_u4_544_wire, CONCAT_u2_u4_571_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_544_wire, CONCAT_u2_u4_571_wire, tmp_var);
      new_bmask_573 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_419_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_418_wire_constant, tmp_var);
      s0_420 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_424_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_423_wire_constant, tmp_var);
      s1_425 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_429_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_428_wire_constant, tmp_var);
      s2_430 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_434_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_433_wire_constant, tmp_var);
      s3_435 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_439_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_438_wire_constant, tmp_var);
      s4_440 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_444_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_443_wire_constant, tmp_var);
      s5_445 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_449_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_448_wire_constant, tmp_var);
      s6_450 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_454_inst
    process(sel_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_368, konst_453_wire_constant, tmp_var);
      s7_455 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_502_inst
    process(lock_val_496) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(lock_val_496, NOT_u8_u8_501_wire_constant, tmp_var);
      EQ_u8_u1_502_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_465_inst
    process(MUX_460_wire, MUX_464_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_460_wire, MUX_464_wire, tmp_var);
      OR_u8_u8_465_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_474_inst
    process(MUX_469_wire, MUX_473_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_469_wire, MUX_473_wire, tmp_var);
      OR_u8_u8_474_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_475_inst
    process(OR_u8_u8_465_wire, OR_u8_u8_474_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_465_wire, OR_u8_u8_474_wire, tmp_var);
      OR_u8_u8_475_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_484_inst
    process(MUX_479_wire, MUX_483_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_479_wire, MUX_483_wire, tmp_var);
      OR_u8_u8_484_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_493_inst
    process(MUX_488_wire, MUX_492_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_488_wire, MUX_492_wire, tmp_var);
      OR_u8_u8_493_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_494_inst
    process(OR_u8_u8_484_wire, OR_u8_u8_493_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_484_wire, OR_u8_u8_493_wire, tmp_var);
      OR_u8_u8_494_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_495_inst
    process(OR_u8_u8_475_wire, OR_u8_u8_494_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_475_wire, OR_u8_u8_494_wire, tmp_var);
      lock_val_496 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_359_call call_stmt_383_call call_stmt_514_call call_stmt_587_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(439 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= call_stmt_359_call_req_0;
      reqL_unguarded(2) <= call_stmt_383_call_req_0;
      reqL_unguarded(1) <= call_stmt_514_call_req_0;
      reqL_unguarded(0) <= call_stmt_587_call_req_0;
      call_stmt_359_call_ack_0 <= ackL_unguarded(3);
      call_stmt_383_call_ack_0 <= ackL_unguarded(2);
      call_stmt_514_call_ack_0 <= ackL_unguarded(1);
      call_stmt_587_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= call_stmt_359_call_req_1;
      reqR_unguarded(2) <= call_stmt_383_call_req_1;
      reqR_unguarded(1) <= call_stmt_514_call_req_1;
      reqR_unguarded(0) <= call_stmt_587_call_req_1;
      call_stmt_359_call_ack_1 <= ackR_unguarded(3);
      call_stmt_383_call_ack_1 <= ackR_unguarded(2);
      call_stmt_514_call_ack_1 <= ackR_unguarded(1);
      call_stmt_587_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_349_wire_constant & type_cast_351_wire_constant & NOT_u8_u8_354_wire_constant & lock_address_pointer_346 & type_cast_357_wire_constant & type_cast_370_wire_constant & type_cast_372_wire_constant & NOT_u8_u8_375_wire_constant & CONCAT_u4_u36_379_wire & type_cast_381_wire_constant & type_cast_504_wire_constant & type_cast_506_wire_constant & NOT_u8_u8_509_wire_constant & lock_address_pointer_346 & type_cast_512_wire_constant & type_cast_575_wire_constant & type_cast_577_wire_constant & new_bmask_573 & CONCAT_u4_u36_582_wire & NOT_u64_u64_585_wire_constant;
      msg_size_plus_lock_359 <= data_out(255 downto 192);
      lock_values_383 <= data_out(191 downto 128);
      err_514 <= data_out(127 downto 64);
      ignore_587 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 440,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 4,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 256,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 4) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(31 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(31 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_1700_start: Boolean;
  signal delay_time_CP_1700_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1390_branch_req_0 : boolean;
  signal phi_stmt_1392_req_1 : boolean;
  signal phi_stmt_1392_req_0 : boolean;
  signal phi_stmt_1392_ack_0 : boolean;
  signal T_1394_buf_req_0 : boolean;
  signal T_1394_buf_ack_0 : boolean;
  signal T_1394_buf_req_1 : boolean;
  signal T_1394_buf_ack_1 : boolean;
  signal nR_1401_1395_buf_req_0 : boolean;
  signal nR_1401_1395_buf_ack_0 : boolean;
  signal nR_1401_1395_buf_req_1 : boolean;
  signal nR_1401_1395_buf_ack_1 : boolean;
  signal do_while_stmt_1390_branch_ack_0 : boolean;
  signal do_while_stmt_1390_branch_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= delay_time_CP_1700_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  delay_time_CP_1700_start <= sample_req;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_1700_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_1700: Block -- control-path 
    signal delay_time_CP_1700_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    delay_time_CP_1700_elements(0) <= delay_time_CP_1700_start;
    delay_time_CP_1700_symbol <= delay_time_CP_1700_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1389/do_while_stmt_1390__entry__
      -- CP-element group 0: 	 branch_block_stmt_1389/branch_block_stmt_1389__entry__
      -- CP-element group 0: 	 branch_block_stmt_1389/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	32 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (8) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1389/assign_stmt_1408__entry__
      -- CP-element group 1: 	 branch_block_stmt_1389/do_while_stmt_1390__exit__
      -- CP-element group 1: 	 branch_block_stmt_1389/$exit
      -- CP-element group 1: 	 branch_block_stmt_1389/assign_stmt_1408__exit__
      -- CP-element group 1: 	 branch_block_stmt_1389/branch_block_stmt_1389__exit__
      -- CP-element group 1: 	 branch_block_stmt_1389/assign_stmt_1408/$entry
      -- CP-element group 1: 	 branch_block_stmt_1389/assign_stmt_1408/$exit
      -- 
    delay_time_CP_1700_elements(1) <= delay_time_CP_1700_elements(32);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1389/do_while_stmt_1390/$entry
      -- CP-element group 2: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390__entry__
      -- 
    delay_time_CP_1700_elements(2) <= delay_time_CP_1700_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	32 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390__exit__
      -- 
    -- Element group delay_time_CP_1700_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_back
      -- 
    -- Element group delay_time_CP_1700_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1389/do_while_stmt_1390/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_taken/$entry
      -- 
    delay_time_CP_1700_elements(5) <= delay_time_CP_1700_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	14 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_body_done
      -- 
    delay_time_CP_1700_elements(6) <= delay_time_CP_1700_elements(14);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/back_edge_to_loop_body
      -- 
    delay_time_CP_1700_elements(7) <= delay_time_CP_1700_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/first_time_through_loop_body
      -- 
    delay_time_CP_1700_elements(8) <= delay_time_CP_1700_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	29 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/loop_body_start
      -- 
    -- Element group delay_time_CP_1700_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	29 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/condition_evaluated
      -- 
    condition_evaluated_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(10), ack => do_while_stmt_1390_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1700_elements(15) & delay_time_CP_1700_elements(29);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1700_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/aggregated_phi_sample_req
      -- 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1700_elements(12) & delay_time_CP_1700_elements(15);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1700_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_sample_start_
      -- 
    delay_time_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1700_elements(9) & delay_time_CP_1700_elements(14);
      gj_delay_time_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1700_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_update_start_
      -- 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1700_elements(9) & delay_time_CP_1700_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1700_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/$exit
      -- CP-element group 14: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_sample_completed__ps
      -- 
    -- Element group delay_time_CP_1700_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_update_completed__ps
      -- 
    -- Element group delay_time_CP_1700_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_loopback_trigger
      -- 
    delay_time_CP_1700_elements(16) <= delay_time_CP_1700_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_loopback_sample_req_ps
      -- 
    phi_stmt_1392_loopback_sample_req_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1392_loopback_sample_req_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(17), ack => phi_stmt_1392_req_1); -- 
    -- Element group delay_time_CP_1700_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_entry_trigger
      -- 
    delay_time_CP_1700_elements(18) <= delay_time_CP_1700_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_entry_sample_req_ps
      -- 
    phi_stmt_1392_entry_sample_req_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1392_entry_sample_req_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(19), ack => phi_stmt_1392_req_0); -- 
    -- Element group delay_time_CP_1700_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/phi_stmt_1392_phi_mux_ack_ps
      -- 
    phi_stmt_1392_phi_mux_ack_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1392_ack_0, ack => delay_time_CP_1700_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Sample/req
      -- 
    req_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(21), ack => T_1394_buf_req_0); -- 
    -- Element group delay_time_CP_1700_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Update/req
      -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(22), ack => T_1394_buf_req_1); -- 
    -- Element group delay_time_CP_1700_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_sample_completed__ps
      -- CP-element group 23: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Sample/ack
      -- 
    ack_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1394_buf_ack_0, ack => delay_time_CP_1700_elements(23)); -- 
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_T_1394_Update/ack
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1394_buf_ack_1, ack => delay_time_CP_1700_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Sample/req
      -- 
    req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(25), ack => nR_1401_1395_buf_req_0); -- 
    -- Element group delay_time_CP_1700_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Update/req
      -- 
    req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1700_elements(26), ack => nR_1401_1395_buf_req_1); -- 
    -- Element group delay_time_CP_1700_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Sample/ack
      -- 
    ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1401_1395_buf_ack_0, ack => delay_time_CP_1700_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/R_nR_1395_Update/ack
      -- 
    ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1401_1395_buf_ack_1, ack => delay_time_CP_1700_elements(28)); -- 
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	10 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1389/do_while_stmt_1390/do_while_stmt_1390_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group delay_time_CP_1700_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => delay_time_CP_1700_elements(9), ack => delay_time_CP_1700_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_exit/$exit
      -- CP-element group 30: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_exit/ack
      -- 
    ack_1790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1390_branch_ack_0, ack => delay_time_CP_1700_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_taken/$exit
      -- CP-element group 31: 	 branch_block_stmt_1389/do_while_stmt_1390/loop_taken/ack
      -- 
    ack_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1390_branch_ack_1, ack => delay_time_CP_1700_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	1 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1389/do_while_stmt_1390/$exit
      -- 
    delay_time_CP_1700_elements(32) <= delay_time_CP_1700_elements(3);
    delay_time_do_while_stmt_1390_terminator_1795: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_1390_terminator_1795", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_1700_elements(6),loop_continue => delay_time_CP_1700_elements(31),loop_terminate => delay_time_CP_1700_elements(30),loop_back => delay_time_CP_1700_elements(4),loop_exit => delay_time_CP_1700_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1392_phi_seq_1785_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_1700_elements(18);
      delay_time_CP_1700_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_1700_elements(23);
      delay_time_CP_1700_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_1700_elements(24);
      delay_time_CP_1700_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_1700_elements(16);
      delay_time_CP_1700_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_1700_elements(27);
      delay_time_CP_1700_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_1700_elements(28);
      delay_time_CP_1700_elements(17) <= phi_mux_reqs(1);
      phi_stmt_1392_phi_seq_1785 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1392_phi_seq_1785") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_1700_elements(11), 
          phi_sample_ack => delay_time_CP_1700_elements(14), 
          phi_update_req => delay_time_CP_1700_elements(13), 
          phi_update_ack => delay_time_CP_1700_elements(15), 
          phi_mux_ack => delay_time_CP_1700_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1727_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_1700_elements(7);
        preds(1)  <= delay_time_CP_1700_elements(8);
        entry_tmerge_1727 : transition_merge -- 
          generic map(name => " entry_tmerge_1727")
          port map (preds => preds, symbol_out => delay_time_CP_1700_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_1392 : std_logic_vector(31 downto 0);
    signal T_1394_buffered : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_1405_wire : std_logic_vector(0 downto 0);
    signal konst_1399_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1404_wire_constant : std_logic_vector(31 downto 0);
    signal nR_1401 : std_logic_vector(31 downto 0);
    signal nR_1401_1395_buffered : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_1399_wire_constant <= "00000000000000000000000000000001";
    konst_1404_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_1392: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= T_1394_buffered & nR_1401_1395_buffered;
      req <= phi_stmt_1392_req_0 & phi_stmt_1392_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1392",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1392_ack_0,
          idata => idata,
          odata => R_1392,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1392
    T_1394_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_1394_buf_req_0;
      T_1394_buf_ack_0<= wack(0);
      rreq(0) <= T_1394_buf_req_1;
      T_1394_buf_ack_1<= rack(0);
      T_1394_buf : InterlockBuffer generic map ( -- 
        name => "T_1394_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_1394_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nR_1401_1395_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_1401_1395_buf_req_0;
      nR_1401_1395_buf_ack_0<= wack(0);
      rreq(0) <= nR_1401_1395_buf_req_1;
      nR_1401_1395_buf_ack_1<= rack(0);
      nR_1401_1395_buf : InterlockBuffer generic map ( -- 
        name => "nR_1401_1395_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_1401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_1401_1395_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1390_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u32_u1_1405_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1390_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1390_branch_req_0,
          ack0 => do_while_stmt_1390_branch_ack_0,
          ack1 => do_while_stmt_1390_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator SUB_u32_u32_1400_inst
    process(R_1392) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_1392, konst_1399_wire_constant, tmp_var);
      nR_1401 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1405_inst
    process(R_1392) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_1392, konst_1404_wire_constant, tmp_var);
      UGT_u32_u1_1405_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    read_index : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal read_index_buffer :  std_logic_vector(31 downto 0);
  signal read_index_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_822_start: Boolean;
  signal getQueueElement_CP_822_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal MUX_727_inst_ack_0 : boolean;
  signal MUX_727_inst_req_0 : boolean;
  signal MUX_727_inst_ack_1 : boolean;
  signal MUX_727_inst_req_1 : boolean;
  signal call_stmt_712_call_ack_1 : boolean;
  signal call_stmt_712_call_req_1 : boolean;
  signal call_stmt_712_call_ack_0 : boolean;
  signal call_stmt_712_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= read_index;
  read_index_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_822_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_822_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_822_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_822_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_822: Block -- control-path 
    signal getQueueElement_CP_822_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_822_elements(0) <= getQueueElement_CP_822_start;
    getQueueElement_CP_822_symbol <= getQueueElement_CP_822_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_complete/$entry
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/$entry
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_sample_start_
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_complete/req
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_update_start_
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_update_start_
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Update/ccr
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Update/$entry
      -- CP-element group 0: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Sample/crr
      -- 
    req_854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_822_elements(0), ack => MUX_727_inst_req_1); -- 
    ccr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_822_elements(0), ack => call_stmt_712_call_req_1); -- 
    crr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_822_elements(0), ack => call_stmt_712_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_sample_completed_
      -- CP-element group 1: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Sample/cra
      -- 
    cra_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_712_call_ack_0, ack => getQueueElement_CP_822_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_start/req
      -- CP-element group 2: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_update_completed_
      -- CP-element group 2: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_start/$entry
      -- CP-element group 2: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_sample_start_
      -- CP-element group 2: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Update/cca
      -- CP-element group 2: 	 assign_stmt_688_to_assign_stmt_728/call_stmt_712_Update/$exit
      -- 
    cca_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_712_call_ack_1, ack => getQueueElement_CP_822_elements(2)); -- 
    req_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_822_elements(2), ack => MUX_727_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_start/ack
      -- CP-element group 3: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_start/$exit
      -- CP-element group 3: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_sample_completed_
      -- 
    ack_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_727_inst_ack_0, ack => getQueueElement_CP_822_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_688_to_assign_stmt_728/$exit
      -- CP-element group 4: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_complete/$exit
      -- CP-element group 4: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_complete/ack
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 assign_stmt_688_to_assign_stmt_728/MUX_727_update_completed_
      -- 
    ack_855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_727_inst_ack_1, ack => getQueueElement_CP_822_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_724_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_696_wire : std_logic_vector(33 downto 0);
    signal NOT_u8_u8_707_wire_constant : std_logic_vector(7 downto 0);
    signal buffer_address_688 : std_logic_vector(35 downto 0);
    signal e0_716 : std_logic_vector(31 downto 0);
    signal e1_720 : std_logic_vector(31 downto 0);
    signal element_pair_712 : std_logic_vector(63 downto 0);
    signal element_pair_address_700 : std_logic_vector(35 downto 0);
    signal konst_723_wire_constant : std_logic_vector(31 downto 0);
    signal slice_693_wire : std_logic_vector(30 downto 0);
    signal type_cast_686_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_695_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_698_wire : std_logic_vector(35 downto 0);
    signal type_cast_702_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_704_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_710_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_707_wire_constant <= "11111111";
    konst_723_wire_constant <= "00000000000000000000000000000000";
    type_cast_686_wire_constant <= "000000000000000000000000000000100000";
    type_cast_695_wire_constant <= "000";
    type_cast_702_wire_constant <= "0";
    type_cast_704_wire_constant <= "1";
    type_cast_710_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    MUX_727_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_727_inst_req_0;
      MUX_727_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_727_inst_req_1;
      MUX_727_inst_ack_1<= update_ack(0);
      MUX_727_inst: SelectSplitProtocol generic map(name => "MUX_727_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => e1_720, y => e0_716, sel => BITSEL_u32_u1_724_wire, z => q_r_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_693_inst
    slice_693_wire <= read_index_buffer(31 downto 1);
    -- flow-through slice operator slice_715_inst
    e0_716 <= element_pair_712(63 downto 32);
    -- flow-through slice operator slice_719_inst
    e1_720 <= element_pair_712(31 downto 0);
    -- interlock type_cast_698_inst
    process(CONCAT_u31_u34_696_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_696_wire(33 downto 0);
      type_cast_698_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_687_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_686_wire_constant, tmp_var);
      buffer_address_688 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_699_inst
    process(buffer_address_688, type_cast_698_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_688, type_cast_698_wire, tmp_var);
      element_pair_address_700 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_724_inst
    process(read_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(read_index_buffer, konst_723_wire_constant, tmp_var);
      BITSEL_u32_u1_724_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_696_inst
    process(slice_693_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_693_wire, type_cast_695_wire_constant, tmp_var);
      CONCAT_u31_u34_696_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_712_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_712_call_req_0;
      call_stmt_712_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_712_call_req_1;
      call_stmt_712_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_702_wire_constant & type_cast_704_wire_constant & NOT_u8_u8_707_wire_constant & element_pair_address_700 & type_cast_710_wire_constant;
      element_pair_712 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueueLength is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    Queue_Length : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueLength;
architecture getQueueLength_arch of getQueueLength is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal Queue_Length_buffer :  std_logic_vector(31 downto 0);
  signal Queue_Length_update_enable: Boolean;
  signal getQueueLength_CP_754_start: Boolean;
  signal getQueueLength_CP_754_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_653_call_req_0 : boolean;
  signal call_stmt_653_call_ack_0 : boolean;
  signal call_stmt_653_call_req_1 : boolean;
  signal call_stmt_653_call_ack_1 : boolean;
  signal slice_656_inst_req_0 : boolean;
  signal slice_656_inst_ack_0 : boolean;
  signal slice_656_inst_req_1 : boolean;
  signal slice_656_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueLength_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueLength_CP_754_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueLength_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= Queue_Length_buffer;
  Queue_Length <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_754_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueLength_CP_754_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_754_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueLength_CP_754: Block -- control-path 
    signal getQueueLength_CP_754_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueLength_CP_754_elements(0) <= getQueueLength_CP_754_start;
    getQueueLength_CP_754_symbol <= getQueueLength_CP_754_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/$entry
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_sample_start_
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_update_start_
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Sample/$entry
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Sample/crr
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Update/$entry
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Update/ccr
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/slice_656_update_start_
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/slice_656_Update/$entry
      -- CP-element group 0: 	 call_stmt_653_to_assign_stmt_657/slice_656_Update/cr
      -- 
    crr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_754_elements(0), ack => call_stmt_653_call_req_0); -- 
    ccr_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_754_elements(0), ack => call_stmt_653_call_req_1); -- 
    cr_786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_754_elements(0), ack => slice_656_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_sample_completed_
      -- CP-element group 1: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Sample/$exit
      -- CP-element group 1: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Sample/cra
      -- 
    cra_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_653_call_ack_0, ack => getQueueLength_CP_754_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_update_completed_
      -- CP-element group 2: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Update/$exit
      -- CP-element group 2: 	 call_stmt_653_to_assign_stmt_657/call_stmt_653_Update/cca
      -- CP-element group 2: 	 call_stmt_653_to_assign_stmt_657/slice_656_sample_start_
      -- CP-element group 2: 	 call_stmt_653_to_assign_stmt_657/slice_656_Sample/$entry
      -- CP-element group 2: 	 call_stmt_653_to_assign_stmt_657/slice_656_Sample/rr
      -- 
    cca_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_653_call_ack_1, ack => getQueueLength_CP_754_elements(2)); -- 
    rr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_754_elements(2), ack => slice_656_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_653_to_assign_stmt_657/slice_656_sample_completed_
      -- CP-element group 3: 	 call_stmt_653_to_assign_stmt_657/slice_656_Sample/$exit
      -- CP-element group 3: 	 call_stmt_653_to_assign_stmt_657/slice_656_Sample/ra
      -- 
    ra_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_656_inst_ack_0, ack => getQueueLength_CP_754_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_653_to_assign_stmt_657/$exit
      -- CP-element group 4: 	 call_stmt_653_to_assign_stmt_657/slice_656_update_completed_
      -- CP-element group 4: 	 call_stmt_653_to_assign_stmt_657/slice_656_Update/$exit
      -- CP-element group 4: 	 call_stmt_653_to_assign_stmt_657/slice_656_Update/ca
      -- 
    ca_787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_656_inst_ack_1, ack => getQueueLength_CP_754_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_649_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_646_wire_constant : std_logic_vector(7 downto 0);
    signal konst_648_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_643_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_651_wire_constant : std_logic_vector(63 downto 0);
    signal wi_and_len_653 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_646_wire_constant <= "11111111";
    konst_648_wire_constant <= "000000000000000000000000000000001000";
    type_cast_641_wire_constant <= "0";
    type_cast_643_wire_constant <= "1";
    type_cast_651_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_656_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_656_inst_req_0;
      slice_656_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_656_inst_req_1;
      slice_656_inst_ack_1<= update_ack(0);
      slice_656_inst: SliceSplitProtocol generic map(name => "slice_656_inst", in_data_width => 64, high_index => 31, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => wi_and_len_653, dout => Queue_Length_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- binary operator ADD_u36_u36_649_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_648_wire_constant, tmp_var);
      ADD_u36_u36_649_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_653_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_653_call_req_0;
      call_stmt_653_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_653_call_req_1;
      call_stmt_653_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_641_wire_constant & type_cast_643_wire_constant & NOT_u8_u8_646_wire_constant & ADD_u36_u36_649_wire & type_cast_651_wire_constant;
      wi_and_len_653 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueLength_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_720_start: Boolean;
  signal getQueuePointers_CP_720_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_609_call_req_0 : boolean;
  signal call_stmt_609_call_ack_0 : boolean;
  signal call_stmt_609_call_req_1 : boolean;
  signal call_stmt_609_call_ack_1 : boolean;
  signal call_stmt_623_call_req_0 : boolean;
  signal call_stmt_623_call_ack_0 : boolean;
  signal call_stmt_623_call_req_1 : boolean;
  signal call_stmt_623_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_720_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_720_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_720_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_720_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_720: Block -- control-path 
    signal getQueuePointers_CP_720_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_720_elements(0) <= getQueuePointers_CP_720_start;
    getQueuePointers_CP_720_symbol <= getQueuePointers_CP_720_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/$entry
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_sample_start_
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_update_start_
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Sample/$entry
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Sample/crr
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Update/$entry
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Update/ccr
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_update_start_
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Update/$entry
      -- CP-element group 0: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Update/ccr
      -- 
    ccr_752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_720_elements(0), ack => call_stmt_623_call_req_1); -- 
    crr_733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_720_elements(0), ack => call_stmt_609_call_req_0); -- 
    ccr_738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_720_elements(0), ack => call_stmt_609_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_sample_completed_
      -- CP-element group 1: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Sample/$exit
      -- CP-element group 1: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Sample/cra
      -- 
    cra_734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_609_call_ack_0, ack => getQueuePointers_CP_720_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_update_completed_
      -- CP-element group 2: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Update/$exit
      -- CP-element group 2: 	 call_stmt_609_to_assign_stmt_631/call_stmt_609_Update/cca
      -- CP-element group 2: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_sample_start_
      -- CP-element group 2: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Sample/$entry
      -- CP-element group 2: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Sample/crr
      -- 
    cca_739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_609_call_ack_1, ack => getQueuePointers_CP_720_elements(2)); -- 
    crr_747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_720_elements(2), ack => call_stmt_623_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_sample_completed_
      -- CP-element group 3: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Sample/$exit
      -- CP-element group 3: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Sample/cra
      -- 
    cra_748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_623_call_ack_0, ack => getQueuePointers_CP_720_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_609_to_assign_stmt_631/$exit
      -- CP-element group 4: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_update_completed_
      -- CP-element group 4: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Update/$exit
      -- CP-element group 4: 	 call_stmt_609_to_assign_stmt_631/call_stmt_623_Update/cca
      -- 
    cca_753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_623_call_ack_1, ack => getQueuePointers_CP_720_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_619_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_604_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_616_wire_constant : std_logic_vector(7 downto 0);
    signal konst_618_wire_constant : std_logic_vector(35 downto 0);
    signal msgs_rp_609 : std_logic_vector(63 downto 0);
    signal type_cast_599_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_601_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_611_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_613_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_621_wire_constant : std_logic_vector(63 downto 0);
    signal wp_len_623 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_604_wire_constant <= "11111111";
    NOT_u8_u8_616_wire_constant <= "11111111";
    konst_618_wire_constant <= "000000000000000000000000000000001000";
    type_cast_599_wire_constant <= "0";
    type_cast_601_wire_constant <= "1";
    type_cast_607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_611_wire_constant <= "0";
    type_cast_613_wire_constant <= "1";
    type_cast_621_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through slice operator slice_626_inst
    rp_buffer <= msgs_rp_609(31 downto 0);
    -- flow-through slice operator slice_630_inst
    wp_buffer <= wp_len_623(63 downto 32);
    -- binary operator ADD_u36_u36_619_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_618_wire_constant, tmp_var);
      ADD_u36_u36_619_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_609_call call_stmt_623_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_609_call_req_0;
      reqL_unguarded(0) <= call_stmt_623_call_req_0;
      call_stmt_609_call_ack_0 <= ackL_unguarded(1);
      call_stmt_623_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_609_call_req_1;
      reqR_unguarded(0) <= call_stmt_623_call_req_1;
      call_stmt_609_call_ack_1 <= ackR_unguarded(1);
      call_stmt_623_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_599_wire_constant & type_cast_601_wire_constant & NOT_u8_u8_604_wire_constant & q_base_address_buffer & type_cast_607_wire_constant & type_cast_611_wire_constant & type_cast_613_wire_constant & NOT_u8_u8_616_wire_constant & ADD_u36_u36_619_wire & type_cast_621_wire_constant;
      msgs_rp_609 <= data_out(127 downto 64);
      wp_len_623 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    total_msgs : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTotalMessages;
architecture getTotalMessages_arch of getTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal total_msgs_update_enable: Boolean;
  signal getTotalMessages_CP_788_start: Boolean;
  signal getTotalMessages_CP_788_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal slice_676_inst_req_1 : boolean;
  signal call_stmt_673_call_ack_0 : boolean;
  signal slice_676_inst_ack_1 : boolean;
  signal slice_676_inst_req_0 : boolean;
  signal call_stmt_673_call_req_0 : boolean;
  signal slice_676_inst_ack_0 : boolean;
  signal call_stmt_673_call_req_1 : boolean;
  signal call_stmt_673_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTotalMessages_CP_788_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= total_msgs_buffer;
  total_msgs <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_788_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTotalMessages_CP_788_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_788_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTotalMessages_CP_788: Block -- control-path 
    signal getTotalMessages_CP_788_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getTotalMessages_CP_788_elements(0) <= getTotalMessages_CP_788_start;
    getTotalMessages_CP_788_symbol <= getTotalMessages_CP_788_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/slice_676_Update/$entry
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/slice_676_Update/cr
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Sample/$entry
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_sample_start_
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_update_start_
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/$entry
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Update/$entry
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Sample/crr
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Update/ccr
      -- CP-element group 0: 	 call_stmt_673_to_assign_stmt_677/slice_676_update_start_
      -- CP-element group 0: 	 $entry
      -- 
    crr_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_788_elements(0), ack => call_stmt_673_call_req_0); -- 
    ccr_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_788_elements(0), ack => call_stmt_673_call_req_1); -- 
    cr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_788_elements(0), ack => slice_676_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Sample/cra
      -- CP-element group 1: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_sample_completed_
      -- CP-element group 1: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Sample/$exit
      -- 
    cra_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_673_call_ack_0, ack => getTotalMessages_CP_788_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_673_to_assign_stmt_677/slice_676_Sample/rr
      -- CP-element group 2: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_update_completed_
      -- CP-element group 2: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Update/$exit
      -- CP-element group 2: 	 call_stmt_673_to_assign_stmt_677/call_stmt_673_Update/cca
      -- CP-element group 2: 	 call_stmt_673_to_assign_stmt_677/slice_676_sample_start_
      -- CP-element group 2: 	 call_stmt_673_to_assign_stmt_677/slice_676_Sample/$entry
      -- 
    cca_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_673_call_ack_1, ack => getTotalMessages_CP_788_elements(2)); -- 
    rr_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_788_elements(2), ack => slice_676_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_673_to_assign_stmt_677/slice_676_Sample/ra
      -- CP-element group 3: 	 call_stmt_673_to_assign_stmt_677/slice_676_sample_completed_
      -- CP-element group 3: 	 call_stmt_673_to_assign_stmt_677/slice_676_Sample/$exit
      -- 
    ra_816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_676_inst_ack_0, ack => getTotalMessages_CP_788_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 call_stmt_673_to_assign_stmt_677/slice_676_Update/ca
      -- CP-element group 4: 	 call_stmt_673_to_assign_stmt_677/slice_676_Update/$exit
      -- CP-element group 4: 	 call_stmt_673_to_assign_stmt_677/$exit
      -- CP-element group 4: 	 call_stmt_673_to_assign_stmt_677/slice_676_update_completed_
      -- CP-element group 4: 	 $exit
      -- 
    ca_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_676_inst_ack_1, ack => getTotalMessages_CP_788_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u8_u8_668_wire_constant : std_logic_vector(7 downto 0);
    signal rdata_673 : std_logic_vector(63 downto 0);
    signal type_cast_663_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_671_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_668_wire_constant <= "11111111";
    type_cast_663_wire_constant <= "0";
    type_cast_665_wire_constant <= "1";
    type_cast_671_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_676_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_676_inst_req_0;
      slice_676_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_676_inst_req_1;
      slice_676_inst_ack_1<= update_ack(0);
      slice_676_inst: SliceSplitProtocol generic map(name => "slice_676_inst", in_data_width => 64, high_index => 63, low_index => 32, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdata_673, dout => total_msgs_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared call operator group (0) : call_stmt_673_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_673_call_req_0;
      call_stmt_673_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_673_call_req_1;
      call_stmt_673_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_663_wire_constant & type_cast_665_wire_constant & NOT_u8_u8_668_wire_constant & q_base_address_buffer & type_cast_671_wire_constant;
      rdata_673 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_index : in  std_logic_vector(5 downto 0);
    pkt_pointer : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_index_buffer :  std_logic_vector(5 downto 0);
  signal queue_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(31 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_3220_start: Boolean;
  signal getTxPacketPointerFromServer_CP_3220_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1858_call_req_0 : boolean;
  signal call_stmt_1858_call_ack_0 : boolean;
  signal call_stmt_1858_call_req_1 : boolean;
  signal call_stmt_1858_call_ack_1 : boolean;
  signal call_stmt_1870_call_req_0 : boolean;
  signal call_stmt_1870_call_ack_0 : boolean;
  signal call_stmt_1870_call_req_1 : boolean;
  signal call_stmt_1870_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= queue_index;
  queue_index_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 7);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= queue_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_3220_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_3220_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_3220_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_3220_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_3220: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_3220_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_3220_elements(0) <= getTxPacketPointerFromServer_CP_3220_start;
    getTxPacketPointerFromServer_CP_3220_symbol <= getTxPacketPointerFromServer_CP_3220_elements(16);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_1848_to_stmt_1875/$entry
      -- 
    getTxPacketPointerFromServer_CP_3220_elements(1) <= getTxPacketPointerFromServer_CP_3220_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_1848_to_stmt_1875/queue_index_update_enable
      -- CP-element group 2: 	 assign_stmt_1848_to_stmt_1875/queue_index_update_enable_out
      -- 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_3220_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3220_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_1848_to_stmt_1875/pkt_pointer_update_enable
      -- CP-element group 3: 	 assign_stmt_1848_to_stmt_1875/pkt_pointer_update_enable_in
      -- 
    getTxPacketPointerFromServer_CP_3220_elements(3) <= getTxPacketPointerFromServer_CP_3220_elements(14);
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_1848_to_stmt_1875/status_update_enable
      -- CP-element group 4: 	 assign_stmt_1848_to_stmt_1875/status_update_enable_in
      -- 
    getTxPacketPointerFromServer_CP_3220_elements(4) <= getTxPacketPointerFromServer_CP_3220_elements(15);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_sample_start_
      -- CP-element group 5: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Sample/crr
      -- 
    crr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_3220_elements(5), ack => call_stmt_1858_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_3220_elements(1) & getTxPacketPointerFromServer_CP_3220_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3220_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_update_start_
      -- CP-element group 6: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Update/$entry
      -- CP-element group 6: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Update/ccr
      -- 
    ccr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_3220_elements(6), ack => call_stmt_1858_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_3220_elements(8) & getTxPacketPointerFromServer_CP_3220_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3220_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_sample_completed_
      -- CP-element group 7: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Sample/cra
      -- 
    cra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1858_call_ack_0, ack => getTxPacketPointerFromServer_CP_3220_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_update_completed_
      -- CP-element group 8: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Update/$exit
      -- CP-element group 8: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1858_Update/cca
      -- 
    cca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1858_call_ack_1, ack => getTxPacketPointerFromServer_CP_3220_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_sample_start_
      -- CP-element group 9: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Sample/crr
      -- 
    crr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_3220_elements(9), ack => call_stmt_1870_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_3220_elements(8) & getTxPacketPointerFromServer_CP_3220_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3220_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_update_start_
      -- CP-element group 10: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Update/$entry
      -- CP-element group 10: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Update/ccr
      -- 
    ccr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_3220_elements(10), ack => call_stmt_1870_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "getTxPacketPointerFromServer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_3220_elements(3) & getTxPacketPointerFromServer_CP_3220_elements(4) & getTxPacketPointerFromServer_CP_3220_elements(12);
      gj_getTxPacketPointerFromServer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_3220_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_sample_completed_
      -- CP-element group 11: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Sample/cra
      -- 
    cra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1870_call_ack_0, ack => getTxPacketPointerFromServer_CP_3220_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_1848_to_stmt_1875/$exit
      -- CP-element group 12: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_update_completed_
      -- CP-element group 12: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Update/$exit
      -- CP-element group 12: 	 assign_stmt_1848_to_stmt_1875/call_stmt_1870_Update/cca
      -- 
    cca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1870_call_ack_1, ack => getTxPacketPointerFromServer_CP_3220_elements(12)); -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_CP_3220_elements(13) <= getTxPacketPointerFromServer_CP_3220_elements(2);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 pkt_pointer_update_enable
      -- 
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 status_update_enable
      -- 
    -- CP-element group 16:  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 $exit
      -- 
    getTxPacketPointerFromServer_CP_3220_elements(16) <= getTxPacketPointerFromServer_CP_3220_elements(12);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_3220_elements(14) <= pkt_pointer_update_enable;
    getTxPacketPointerFromServer_CP_3220_elements(15) <= status_update_enable;
    -- hookup: output from control-path 
    queue_index_update_enable <= getTxPacketPointerFromServer_CP_3220_elements(13);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1846_wire : std_logic_vector(5 downto 0);
    signal NOT_u4_u4_1853_wire_constant : std_logic_vector(3 downto 0);
    signal R_TX_QUEUES_REG_START_OFFSET_1845_wire_constant : std_logic_vector(5 downto 0);
    signal register_index_1848 : std_logic_vector(5 downto 0);
    signal tx_queue_pointer_32_1858 : std_logic_vector(31 downto 0);
    signal tx_queue_pointer_36_1864 : std_logic_vector(35 downto 0);
    signal type_cast_1850_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1856_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1861_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1866_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1853_wire_constant <= "1111";
    R_TX_QUEUES_REG_START_OFFSET_1845_wire_constant <= "001010";
    type_cast_1850_wire_constant <= "1";
    type_cast_1856_wire_constant <= "00000000000000000000000000000000";
    type_cast_1861_wire_constant <= "0000";
    type_cast_1866_wire_constant <= "1";
    -- interlock type_cast_1847_inst
    process(ADD_u6_u6_1846_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1846_wire(5 downto 0);
      register_index_1848 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u6_u6_1846_inst
    process(queue_index_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(queue_index_buffer, R_TX_QUEUES_REG_START_OFFSET_1845_wire_constant, tmp_var);
      ADD_u6_u6_1846_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1863_inst
    process(type_cast_1861_wire_constant, tx_queue_pointer_32_1858) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1861_wire_constant, tx_queue_pointer_32_1858, tmp_var);
      tx_queue_pointer_36_1864 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1858_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1858_call_req_0;
      call_stmt_1858_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1858_call_req_1;
      call_stmt_1858_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1850_wire_constant & NOT_u4_u4_1853_wire_constant & register_index_1848 & type_cast_1856_wire_constant;
      tx_queue_pointer_32_1858 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1870_call 
    popFromQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1870_call_req_0;
      call_stmt_1870_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1870_call_req_1;
      call_stmt_1870_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_1_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1866_wire_constant & tx_queue_pointer_36_1864;
      pkt_pointer_buffer <= data_out(32 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(54 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_1432_start: Boolean;
  signal loadBuffer_CP_1432_symbol: Boolean;
  -- volatile/operator module components. 
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(10 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position_out : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(10 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1198_call_req_0 : boolean;
  signal call_stmt_1198_call_ack_0 : boolean;
  signal call_stmt_1198_call_req_1 : boolean;
  signal call_stmt_1198_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_ack_1 : boolean;
  signal call_stmt_1207_call_req_0 : boolean;
  signal call_stmt_1207_call_ack_0 : boolean;
  signal call_stmt_1207_call_req_1 : boolean;
  signal call_stmt_1207_call_ack_1 : boolean;
  signal W_bad_packet_identifier_1210_delayed_8_0_1208_inst_req_0 : boolean;
  signal W_bad_packet_identifier_1210_delayed_8_0_1208_inst_ack_0 : boolean;
  signal W_bad_packet_identifier_1210_delayed_8_0_1208_inst_req_1 : boolean;
  signal W_bad_packet_identifier_1210_delayed_8_0_1208_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_ack_1 : boolean;
  signal call_stmt_1218_call_req_0 : boolean;
  signal call_stmt_1218_call_ack_0 : boolean;
  signal call_stmt_1218_call_req_1 : boolean;
  signal call_stmt_1218_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 31);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_1432_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1432_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_1432_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1432_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_1432: Block -- control-path 
    signal loadBuffer_CP_1432_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_1432_elements(0) <= loadBuffer_CP_1432_start;
    loadBuffer_CP_1432_symbol <= loadBuffer_CP_1432_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	20 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1198_to_call_stmt_1218/$entry
      -- 
    loadBuffer_CP_1432_elements(1) <= loadBuffer_CP_1432_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	22 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1198_to_call_stmt_1218/rx_buffer_pointer_update_enable
      -- CP-element group 2: 	 call_stmt_1198_to_call_stmt_1218/rx_buffer_pointer_update_enable_out
      -- 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(6) & loadBuffer_CP_1432_elements(10) & loadBuffer_CP_1432_elements(22);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	29 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1198_to_call_stmt_1218/bad_packet_identifier_update_enable
      -- CP-element group 3: 	 call_stmt_1198_to_call_stmt_1218/bad_packet_identifier_update_enable_in
      -- 
    loadBuffer_CP_1432_elements(3) <= loadBuffer_CP_1432_elements(29);
    -- CP-element group 4:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	27 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_sample_start_
      -- CP-element group 4: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Sample/crr
      -- 
    crr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(4), ack => call_stmt_1198_call_req_0); -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(1) & loadBuffer_CP_1432_elements(6) & loadBuffer_CP_1432_elements(27);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	14 
    -- CP-element group 5: 	27 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_update_start_
      -- CP-element group 5: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Update/$entry
      -- CP-element group 5: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Update/ccr
      -- 
    ccr_1454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(5), ack => call_stmt_1198_call_req_1); -- 
    loadBuffer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(7) & loadBuffer_CP_1432_elements(14) & loadBuffer_CP_1432_elements(27);
      gj_loadBuffer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: 	4 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_sample_completed_
      -- CP-element group 6: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Sample/$exit
      -- CP-element group 6: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Sample/cra
      -- 
    cra_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1198_call_ack_0, ack => loadBuffer_CP_1432_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_update_completed_
      -- CP-element group 7: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Update/$exit
      -- CP-element group 7: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1198_Update/cca
      -- 
    cca_1455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1198_call_ack_1, ack => loadBuffer_CP_1432_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_sample_start_
      -- CP-element group 8: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Sample/req
      -- 
    req_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(8), ack => W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_req_0); -- 
    loadBuffer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(1) & loadBuffer_CP_1432_elements(10);
      gj_loadBuffer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_update_start_
      -- CP-element group 9: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Update/$entry
      -- CP-element group 9: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Update/req
      -- 
    req_1468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(9), ack => W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_req_1); -- 
    loadBuffer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(11) & loadBuffer_CP_1432_elements(14);
      gj_loadBuffer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_sample_completed_
      -- CP-element group 10: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Sample/$exit
      -- CP-element group 10: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Sample/ack
      -- 
    ack_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_ack_0, ack => loadBuffer_CP_1432_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_update_completed_
      -- CP-element group 11: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Update/$exit
      -- CP-element group 11: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1201_Update/ack
      -- 
    ack_1469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_ack_1, ack => loadBuffer_CP_1432_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_sample_start_
      -- CP-element group 12: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Sample/$entry
      -- CP-element group 12: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Sample/crr
      -- 
    crr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(12), ack => call_stmt_1207_call_req_0); -- 
    loadBuffer_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(7) & loadBuffer_CP_1432_elements(11) & loadBuffer_CP_1432_elements(14);
      gj_loadBuffer_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	26 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_update_start_
      -- CP-element group 13: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Update/$entry
      -- CP-element group 13: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Update/ccr
      -- 
    ccr_1482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(13), ack => call_stmt_1207_call_req_1); -- 
    loadBuffer_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(3) & loadBuffer_CP_1432_elements(15) & loadBuffer_CP_1432_elements(18) & loadBuffer_CP_1432_elements(26);
      gj_loadBuffer_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	5 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_sample_completed_
      -- CP-element group 14: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Sample/$exit
      -- CP-element group 14: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Sample/cra
      -- 
    cra_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1207_call_ack_0, ack => loadBuffer_CP_1432_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	24 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_update_completed_
      -- CP-element group 15: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Update/$exit
      -- CP-element group 15: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1207_Update/cca
      -- 
    cca_1483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1207_call_ack_1, ack => loadBuffer_CP_1432_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_sample_start_
      -- CP-element group 16: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Sample/$entry
      -- CP-element group 16: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Sample/req
      -- 
    req_1491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(16), ack => W_bad_packet_identifier_1210_delayed_8_0_1208_inst_req_0); -- 
    loadBuffer_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(15) & loadBuffer_CP_1432_elements(18);
      gj_loadBuffer_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	26 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_update_start_
      -- CP-element group 17: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Update/$entry
      -- CP-element group 17: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Update/req
      -- 
    req_1496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(17), ack => W_bad_packet_identifier_1210_delayed_8_0_1208_inst_req_1); -- 
    loadBuffer_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(19) & loadBuffer_CP_1432_elements(26);
      gj_loadBuffer_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_sample_completed_
      -- CP-element group 18: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Sample/ack
      -- 
    ack_1492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1210_delayed_8_0_1208_inst_ack_0, ack => loadBuffer_CP_1432_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_update_completed_
      -- CP-element group 19: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Update/$exit
      -- CP-element group 19: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1210_Update/ack
      -- 
    ack_1497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1210_delayed_8_0_1208_inst_ack_1, ack => loadBuffer_CP_1432_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	1 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_sample_start_
      -- CP-element group 20: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Sample/$entry
      -- CP-element group 20: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Sample/req
      -- 
    req_1505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(20), ack => W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_req_0); -- 
    loadBuffer_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(1) & loadBuffer_CP_1432_elements(22);
      gj_loadBuffer_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_update_start_
      -- CP-element group 21: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Update/$entry
      -- CP-element group 21: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Update/req
      -- 
    req_1510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(21), ack => W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_req_1); -- 
    loadBuffer_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(23) & loadBuffer_CP_1432_elements(26);
      gj_loadBuffer_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_sample_completed_
      -- CP-element group 22: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Sample/$exit
      -- CP-element group 22: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Sample/ack
      -- 
    ack_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_ack_0, ack => loadBuffer_CP_1432_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_update_completed_
      -- CP-element group 23: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Update/$exit
      -- CP-element group 23: 	 call_stmt_1198_to_call_stmt_1218/assign_stmt_1213_Update/ack
      -- 
    ack_1511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_ack_1, ack => loadBuffer_CP_1432_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_sample_start_
      -- CP-element group 24: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Sample/$entry
      -- CP-element group 24: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Sample/crr
      -- 
    crr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(24), ack => call_stmt_1218_call_req_0); -- 
    loadBuffer_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1432_elements(15) & loadBuffer_CP_1432_elements(19) & loadBuffer_CP_1432_elements(23) & loadBuffer_CP_1432_elements(26);
      gj_loadBuffer_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_update_start_
      -- CP-element group 25: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Update/$entry
      -- CP-element group 25: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Update/ccr
      -- 
    ccr_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1432_elements(25), ack => call_stmt_1218_call_req_1); -- 
    loadBuffer_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_1432_elements(27);
      gj_loadBuffer_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1432_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: 	17 
    -- CP-element group 26: 	21 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_sample_completed_
      -- CP-element group 26: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Sample/$exit
      -- CP-element group 26: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Sample/cra
      -- 
    cra_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1218_call_ack_0, ack => loadBuffer_CP_1432_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	4 
    -- CP-element group 27: 	5 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 call_stmt_1198_to_call_stmt_1218/$exit
      -- CP-element group 27: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_update_completed_
      -- CP-element group 27: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Update/$exit
      -- CP-element group 27: 	 call_stmt_1198_to_call_stmt_1218/call_stmt_1218_Update/cca
      -- 
    cca_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1218_call_ack_1, ack => loadBuffer_CP_1432_elements(27)); -- 
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 rx_buffer_pointer_update_enable
      -- 
    loadBuffer_CP_1432_elements(28) <= loadBuffer_CP_1432_elements(2);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	3 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 bad_packet_identifier_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    loadBuffer_CP_1432_elements(30) <= loadBuffer_CP_1432_elements(27);
    --  hookup: inputs to control-path 
    loadBuffer_CP_1432_elements(29) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_1432_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal bad_packet_identifier_1210_delayed_8_0_1210 : std_logic_vector(0 downto 0);
    signal last_keep_1207 : std_logic_vector(7 downto 0);
    signal new_buf_pointer_1198 : std_logic_vector(35 downto 0);
    signal packet_size_1207 : std_logic_vector(10 downto 0);
    signal rx_buffer_pointer_1204_delayed_4_0_1201 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_1211_delayed_8_0_1213 : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    W_bad_packet_identifier_1210_delayed_8_0_1208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bad_packet_identifier_1210_delayed_8_0_1208_inst_req_0;
      W_bad_packet_identifier_1210_delayed_8_0_1208_inst_ack_0<= wack(0);
      rreq(0) <= W_bad_packet_identifier_1210_delayed_8_0_1208_inst_req_1;
      W_bad_packet_identifier_1210_delayed_8_0_1208_inst_ack_1<= rack(0);
      W_bad_packet_identifier_1210_delayed_8_0_1208_inst : InterlockBuffer generic map ( -- 
        name => "W_bad_packet_identifier_1210_delayed_8_0_1208_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bad_packet_identifier_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bad_packet_identifier_1210_delayed_8_0_1210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_req_0;
      W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_req_1;
      W_rx_buffer_pointer_1204_delayed_4_0_1199_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1204_delayed_4_0_1199_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1204_delayed_4_0_1199_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1204_delayed_4_0_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_req_0;
      W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_req_1;
      W_rx_buffer_pointer_1211_delayed_8_0_1211_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1211_delayed_8_0_1211_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1211_delayed_8_0_1211_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1211_delayed_8_0_1213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared call operator group (0) : call_stmt_1198_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1198_call_req_0;
      call_stmt_1198_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1198_call_req_1;
      call_stmt_1198_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer;
      new_buf_pointer_1198 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(35 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(35 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1207_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(19 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1207_call_req_0;
      call_stmt_1207_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1207_call_req_1;
      call_stmt_1207_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_1204_delayed_4_0_1201 & new_buf_pointer_1198;
      packet_size_1207 <= data_out(19 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_1207 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(71 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 20,
          owidth => 20,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(19 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1218_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(54 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1218_call_req_0;
      call_stmt_1218_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1218_call_req_1;
      call_stmt_1218_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_1210_delayed_8_0_1210(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_1211_delayed_8_0_1213 & packet_size_1207 & last_keep_1207;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 55,
        owidth => 55,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(54 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1932_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1940_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1896_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1914_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1905_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1911_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1922_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1929_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1938_wire : std_logic_vector(0 downto 0);
    signal MUX_1908_wire : std_logic_vector(1 downto 0);
    signal MUX_1918_wire : std_logic_vector(1 downto 0);
    signal MUX_1925_wire : std_logic_vector(1 downto 0);
    signal MUX_1935_wire : std_logic_vector(1 downto 0);
    signal MUX_1943_wire : std_logic_vector(1 downto 0);
    signal NEQ_u2_u1_1899_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1931_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1915_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_1919_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_1926_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_1944_wire : std_logic_vector(1 downto 0);
    signal R_S0_1904_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1916_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1941_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1906_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1921_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1898_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1923_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1928_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1933_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1937_wire_constant : std_logic_vector(1 downto 0);
    signal R_S3_1910_wire_constant : std_logic_vector(1 downto 0);
    signal go_to_s0_1901 : std_logic_vector(0 downto 0);
    signal konst_1890_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1895_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1907_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1913_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1917_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1924_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1934_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1942_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_1892 : std_logic_vector(0 downto 0);
    signal tlast_1887 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_1904_wire_constant <= "00";
    R_S0_1916_wire_constant <= "00";
    R_S0_1941_wire_constant <= "00";
    R_S1_1906_wire_constant <= "01";
    R_S1_1921_wire_constant <= "01";
    R_S2_1898_wire_constant <= "10";
    R_S2_1923_wire_constant <= "10";
    R_S2_1928_wire_constant <= "10";
    R_S2_1933_wire_constant <= "10";
    R_S2_1937_wire_constant <= "10";
    R_S3_1910_wire_constant <= "11";
    konst_1890_wire_constant <= "1";
    konst_1895_wire_constant <= "1";
    konst_1907_wire_constant <= "00";
    konst_1913_wire_constant <= "1";
    konst_1917_wire_constant <= "00";
    konst_1924_wire_constant <= "00";
    konst_1934_wire_constant <= "00";
    konst_1942_wire_constant <= "00";
    -- flow-through select operator MUX_1908_inst
    MUX_1908_wire <= R_S1_1906_wire_constant when (EQ_u2_u1_1905_wire(0) /=  '0') else konst_1907_wire_constant;
    -- flow-through select operator MUX_1918_inst
    MUX_1918_wire <= R_S0_1916_wire_constant when (OR_u1_u1_1915_wire(0) /=  '0') else konst_1917_wire_constant;
    -- flow-through select operator MUX_1925_inst
    MUX_1925_wire <= R_S2_1923_wire_constant when (EQ_u2_u1_1922_wire(0) /=  '0') else konst_1924_wire_constant;
    -- flow-through select operator MUX_1935_inst
    MUX_1935_wire <= R_S2_1933_wire_constant when (AND_u1_u1_1932_wire(0) /=  '0') else konst_1934_wire_constant;
    -- flow-through select operator MUX_1943_inst
    MUX_1943_wire <= R_S0_1941_wire_constant when (AND_u1_u1_1940_wire(0) /=  '0') else konst_1942_wire_constant;
    -- flow-through slice operator slice_1886_inst
    tlast_1887 <= RX_buffer(72 downto 72);
    -- binary operator AND_u1_u1_1900_inst
    process(EQ_u1_u1_1896_wire, NEQ_u2_u1_1899_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_1896_wire, NEQ_u2_u1_1899_wire, tmp_var);
      go_to_s0_1901 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1932_inst
    process(EQ_u2_u1_1929_wire, NOT_u1_u1_1931_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1929_wire, NOT_u1_u1_1931_wire, tmp_var);
      AND_u1_u1_1932_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1940_inst
    process(EQ_u2_u1_1938_wire, last_word_1892) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1938_wire, last_word_1892, tmp_var);
      AND_u1_u1_1940_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1891_inst
    process(tlast_1887) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_1887, konst_1890_wire_constant, tmp_var);
      last_word_1892 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1896_inst
    process(last_word_1892) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_word_1892, konst_1895_wire_constant, tmp_var);
      EQ_u1_u1_1896_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1914_inst
    process(go_to_s0_1901) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(go_to_s0_1901, konst_1913_wire_constant, tmp_var);
      EQ_u1_u1_1914_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1905_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_1904_wire_constant, tmp_var);
      EQ_u2_u1_1905_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1911_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S3_1910_wire_constant, tmp_var);
      EQ_u2_u1_1911_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1922_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_1921_wire_constant, tmp_var);
      EQ_u2_u1_1922_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1929_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1928_wire_constant, tmp_var);
      EQ_u2_u1_1929_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1938_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1937_wire_constant, tmp_var);
      EQ_u2_u1_1938_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u2_u1_1899_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSTATE_buffer, R_S2_1898_wire_constant, tmp_var);
      NEQ_u2_u1_1899_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1931_inst
    process(last_word_1892) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_1892, tmp_var);
      NOT_u1_u1_1931_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1915_inst
    process(EQ_u2_u1_1911_wire, EQ_u1_u1_1914_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_1911_wire, EQ_u1_u1_1914_wire, tmp_var);
      OR_u1_u1_1915_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1919_inst
    process(MUX_1908_wire, MUX_1918_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1908_wire, MUX_1918_wire, tmp_var);
      OR_u2_u2_1919_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1926_inst
    process(OR_u2_u2_1919_wire, MUX_1925_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_1919_wire, MUX_1925_wire, tmp_var);
      OR_u2_u2_1926_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1944_inst
    process(MUX_1935_wire, MUX_1943_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1935_wire, MUX_1943_wire, tmp_var);
      OR_u2_u2_1944_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1945_inst
    process(OR_u2_u2_1926_wire, OR_u2_u2_1944_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_1926_wire, OR_u2_u2_1944_wire, tmp_var);
      nLSTATE_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(1 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(1 downto 0);
    AccessRegister_call_data : out  std_logic_vector(85 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(1 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(1 downto 0);
    AccessRegister_return_data : in   std_logic_vector(63 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_3269_start: Boolean;
  signal nicRxFromMacDaemon_CP_3269_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component nextLSTATE_Volatile is -- 
    port ( -- 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal WPIPE_nic_rx_to_packet_2023_inst_ack_0 : boolean;
  signal MUX_2021_inst_req_0 : boolean;
  signal npkt_cnt_2039_1991_buf_req_1 : boolean;
  signal npkt_cnt_2039_1991_buf_ack_0 : boolean;
  signal call_stmt_1979_call_ack_1 : boolean;
  signal nLSTATE_2001_1984_buf_ack_1 : boolean;
  signal call_stmt_2049_call_req_0 : boolean;
  signal npkt_cnt_2039_1991_buf_req_0 : boolean;
  signal call_stmt_1961_call_req_1 : boolean;
  signal call_stmt_1979_call_req_0 : boolean;
  signal MUX_2021_inst_ack_0 : boolean;
  signal call_stmt_2049_call_ack_0 : boolean;
  signal npkt_cnt_2039_1991_buf_ack_1 : boolean;
  signal phi_stmt_1982_req_0 : boolean;
  signal if_stmt_1962_branch_req_0 : boolean;
  signal phi_stmt_1989_req_0 : boolean;
  signal do_while_stmt_1980_branch_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_2012_inst_ack_1 : boolean;
  signal MUX_2021_inst_req_1 : boolean;
  signal MUX_2021_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_packet_2023_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_packet_2023_inst_ack_1 : boolean;
  signal call_stmt_2049_call_req_1 : boolean;
  signal if_stmt_1962_branch_ack_1 : boolean;
  signal call_stmt_2049_call_ack_1 : boolean;
  signal phi_stmt_1989_req_1 : boolean;
  signal nLSTATE_2001_1984_buf_req_1 : boolean;
  signal do_while_stmt_1980_branch_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_1988_inst_req_0 : boolean;
  signal if_stmt_1962_branch_ack_0 : boolean;
  signal call_stmt_1979_call_req_1 : boolean;
  signal phi_stmt_1982_req_1 : boolean;
  signal WPIPE_nic_rx_to_header_2012_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1988_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_2012_inst_ack_0 : boolean;
  signal call_stmt_1961_call_req_0 : boolean;
  signal phi_stmt_1982_ack_0 : boolean;
  signal call_stmt_1961_call_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_1988_inst_req_1 : boolean;
  signal phi_stmt_1989_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_2012_inst_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_1988_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_packet_2023_inst_req_0 : boolean;
  signal call_stmt_1961_call_ack_1 : boolean;
  signal nLSTATE_2001_1984_buf_ack_0 : boolean;
  signal do_while_stmt_1980_branch_req_0 : boolean;
  signal nLSTATE_2001_1984_buf_req_0 : boolean;
  signal call_stmt_1979_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_3269_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_3269_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_3269_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_3269_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_3269: Block -- control-path 
    signal nicRxFromMacDaemon_CP_3269_elements: BooleanArray(82 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_3269_elements(0) <= nicRxFromMacDaemon_CP_3269_start;
    nicRxFromMacDaemon_CP_3269_symbol <= nicRxFromMacDaemon_CP_3269_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	82 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1949/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1949/merge_stmt_1951_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1949/branch_block_stmt_1949__entry__
      -- CP-element group 0: 	 branch_block_stmt_1949/merge_stmt_1951__entry__
      -- CP-element group 0: 	 branch_block_stmt_1949/merge_stmt_1951__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1949/merge_stmt_1951__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1949/$exit
      -- CP-element group 1: 	 branch_block_stmt_1949/branch_block_stmt_1949__exit__
      -- CP-element group 1: 	 $exit
      -- 
    nicRxFromMacDaemon_CP_3269_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	81 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	82 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_1949/disable_loopback
      -- CP-element group 2: 	 branch_block_stmt_1949/do_while_stmt_1980__exit__
      -- CP-element group 2: 	 branch_block_stmt_1949/disable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1949/disable_loopback_PhiReq/$exit
      -- 
    nicRxFromMacDaemon_CP_3269_elements(2) <= nicRxFromMacDaemon_CP_3269_elements(81);
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	82 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Sample/cra
      -- 
    cra_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1961_call_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	82 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (49) 
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1949/call_stmt_1961__exit__
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_1949/NOT_u1_u1_1966_place
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Sample/ack
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_else_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Sample/req
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/call_stmt_1961/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962__entry__
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Update/req
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Update/ack
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/BITSEL_u32_u1_1965_inputs/RPIPE_CONTROL_REGISTER_1963/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1949/if_stmt_1962_eval_test/NOT_u1_u1_1966/BITSEL_u32_u1_1965/SplitProtocol/Update/$exit
      -- 
    cca_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1961_call_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(4)); -- 
    branch_req_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(4), ack => if_stmt_1962_branch_req_0); -- 
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	82 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1949/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1949/not_enabled_yet_loopback_PhiReq/$exit
      -- CP-element group 5: 	 branch_block_stmt_1949/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1949/if_stmt_1962_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1949/if_stmt_1962_if_link/if_choice_transition
      -- 
    if_choice_transition_3365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1962_branch_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(5)); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1949/if_stmt_1962_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1949/if_stmt_1962_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/$entry
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Update/ccr
      -- CP-element group 6: 	 branch_block_stmt_1949/if_stmt_1962__exit__
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979__entry__
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Sample/$entry
      -- 
    else_choice_transition_3369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1962_branch_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(6)); -- 
    crr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(6), ack => call_stmt_1979_call_req_0); -- 
    ccr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(6), ack => call_stmt_1979_call_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Sample/cra
      -- 
    cra_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1979_call_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Update/cca
      -- CP-element group 8: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1949/call_stmt_1979/$exit
      -- CP-element group 8: 	 branch_block_stmt_1949/call_stmt_1979__exit__
      -- CP-element group 8: 	 branch_block_stmt_1949/do_while_stmt_1980__entry__
      -- CP-element group 8: 	 branch_block_stmt_1949/call_stmt_1979/call_stmt_1979_update_completed_
      -- 
    cca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1979_call_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(8)); -- 
    -- CP-element group 9:  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980__entry__
      -- CP-element group 9: 	 branch_block_stmt_1949/do_while_stmt_1980/$entry
      -- 
    nicRxFromMacDaemon_CP_3269_elements(9) <= nicRxFromMacDaemon_CP_3269_elements(8);
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	81 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980__exit__
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(10) is bound as output of CP function.
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_back
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(11) is bound as output of CP function.
    -- CP-element group 12:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	80 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1949/do_while_stmt_1980/condition_done
      -- CP-element group 12: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_exit/$entry
      -- CP-element group 12: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_taken/$entry
      -- 
    nicRxFromMacDaemon_CP_3269_elements(12) <= nicRxFromMacDaemon_CP_3269_elements(17);
    -- CP-element group 13:  branch  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	78 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_body_done
      -- 
    nicRxFromMacDaemon_CP_3269_elements(13) <= nicRxFromMacDaemon_CP_3269_elements(78);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	26 
    -- CP-element group 14: 	50 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/back_edge_to_loop_body
      -- 
    nicRxFromMacDaemon_CP_3269_elements(14) <= nicRxFromMacDaemon_CP_3269_elements(11);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	52 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/first_time_through_loop_body
      -- 
    nicRxFromMacDaemon_CP_3269_elements(15) <= nicRxFromMacDaemon_CP_3269_elements(9);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	22 
    -- CP-element group 16: 	23 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	44 
    -- CP-element group 16: 	45 
    -- CP-element group 16: 	77 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1986_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/$entry
      -- CP-element group 16: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/loop_body_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(16) is bound as output of CP function.
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	77 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/condition_evaluated
      -- 
    condition_evaluated_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(17), ack => do_while_stmt_1980_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(21) & nicRxFromMacDaemon_CP_3269_elements(77);
      gj_nicRxFromMacDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	22 
    -- CP-element group 18: 	44 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	40 
    -- CP-element group 18: 	46 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_sample_start__ps
      -- CP-element group 18: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/aggregated_phi_sample_req
      -- 
    nicRxFromMacDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(16) & nicRxFromMacDaemon_CP_3269_elements(22) & nicRxFromMacDaemon_CP_3269_elements(44) & nicRxFromMacDaemon_CP_3269_elements(21);
      gj_nicRxFromMacDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	47 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	78 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	44 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1986_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/aggregated_phi_sample_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(24) & nicRxFromMacDaemon_CP_3269_elements(42) & nicRxFromMacDaemon_CP_3269_elements(47);
      gj_nicRxFromMacDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: 	39 
    -- CP-element group 20: 	45 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	41 
    -- CP-element group 20: 	48 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/aggregated_phi_update_req
      -- CP-element group 20: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_update_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(23) & nicRxFromMacDaemon_CP_3269_elements(39) & nicRxFromMacDaemon_CP_3269_elements(45);
      gj_nicRxFromMacDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	49 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/aggregated_phi_update_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(25) & nicRxFromMacDaemon_CP_3269_elements(43) & nicRxFromMacDaemon_CP_3269_elements(49);
      gj_nicRxFromMacDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(16) & nicRxFromMacDaemon_CP_3269_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	68 
    -- CP-element group 23: 	75 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(16) & nicRxFromMacDaemon_CP_3269_elements(25) & nicRxFromMacDaemon_CP_3269_elements(65) & nicRxFromMacDaemon_CP_3269_elements(68) & nicRxFromMacDaemon_CP_3269_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	21 
    -- CP-element group 25: 	63 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	73 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_update_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_3269_elements(26) <= nicRxFromMacDaemon_CP_3269_elements(14);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_loopback_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_loopback_sample_req_ps
      -- 
    phi_stmt_1982_loopback_sample_req_3417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1982_loopback_sample_req_3417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(27), ack => phi_stmt_1982_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_3269_elements(28) <= nicRxFromMacDaemon_CP_3269_elements(15);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_entry_sample_req
      -- CP-element group 29: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_entry_sample_req_ps
      -- 
    phi_stmt_1982_entry_sample_req_3420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1982_entry_sample_req_3420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(29), ack => phi_stmt_1982_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_phi_mux_ack
      -- CP-element group 30: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1982_phi_mux_ack_ps
      -- 
    phi_stmt_1982_phi_mux_ack_3423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1982_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Sample/req
      -- CP-element group 31: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Sample/$entry
      -- 
    req_3436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(31), ack => nLSTATE_2001_1984_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Update/req
      -- CP-element group 32: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_update_start_
      -- 
    req_3441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(32), ack => nLSTATE_2001_1984_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_sample_completed_
      -- 
    ack_3437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_2001_1984_buf_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_nLSTATE_1984_update_completed_
      -- 
    ack_3442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_2001_1984_buf_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_update_start_
      -- CP-element group 36: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_update_start__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_3269_elements(37) <= nicRxFromMacDaemon_CP_3269_elements(38);
    -- CP-element group 38:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	37 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_S0_1985_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_3269_elements(36), ack => nicRxFromMacDaemon_CP_3269_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	65 
    -- CP-element group 39: 	71 
    -- CP-element group 39: 	75 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	20 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1986_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(16) & nicRxFromMacDaemon_CP_3269_elements(65) & nicRxFromMacDaemon_CP_3269_elements(71) & nicRxFromMacDaemon_CP_3269_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	18 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	43 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Sample/rr
      -- 
    rr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(40), ack => RPIPE_mac_to_nic_data_1988_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(18) & nicRxFromMacDaemon_CP_3269_elements(43);
      gj_nicRxFromMacDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	20 
    -- CP-element group 41: 	42 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Update/cr
      -- 
    cr_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(41), ack => RPIPE_mac_to_nic_data_1988_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(20) & nicRxFromMacDaemon_CP_3269_elements(42);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: 	41 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Sample/ra
      -- 
    ra_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1988_inst_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	21 
    -- CP-element group 43: 	63 
    -- CP-element group 43: 	70 
    -- CP-element group 43: 	73 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	40 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1986_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/RPIPE_mac_to_nic_data_1988_Update/ca
      -- 
    ca_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1988_inst_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(43)); -- 
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	16 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	19 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	18 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(16) & nicRxFromMacDaemon_CP_3269_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	16 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	49 
    -- CP-element group 45: 	75 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	20 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(16) & nicRxFromMacDaemon_CP_3269_elements(49) & nicRxFromMacDaemon_CP_3269_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	18 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_sample_start__ps
      -- 
    nicRxFromMacDaemon_CP_3269_elements(46) <= nicRxFromMacDaemon_CP_3269_elements(18);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	19 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(47) is bound as output of CP function.
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	20 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_update_start__ps
      -- 
    nicRxFromMacDaemon_CP_3269_elements(48) <= nicRxFromMacDaemon_CP_3269_elements(20);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	21 
    -- CP-element group 49: 	73 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	45 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_update_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	14 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_3269_elements(50) <= nicRxFromMacDaemon_CP_3269_elements(14);
    -- CP-element group 51:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_loopback_sample_req
      -- CP-element group 51: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_loopback_sample_req_ps
      -- 
    phi_stmt_1989_loopback_sample_req_3479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1989_loopback_sample_req_3479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(51), ack => phi_stmt_1989_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	15 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_3269_elements(52) <= nicRxFromMacDaemon_CP_3269_elements(15);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_entry_sample_req
      -- CP-element group 53: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_entry_sample_req_ps
      -- 
    phi_stmt_1989_entry_sample_req_3482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1989_entry_sample_req_3482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(53), ack => phi_stmt_1989_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_phi_mux_ack
      -- CP-element group 54: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/phi_stmt_1989_phi_mux_ack_ps
      -- 
    phi_stmt_1989_phi_mux_ack_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1989_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Sample/req
      -- CP-element group 55: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_sample_start_
      -- 
    req_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(55), ack => npkt_cnt_2039_1991_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Update/req
      -- CP-element group 56: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_update_start_
      -- 
    req_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(56), ack => npkt_cnt_2039_1991_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_sample_completed_
      -- 
    ack_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_2039_1991_buf_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/R_npkt_cnt_1991_update_completed__ps
      -- 
    ack_3504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_2039_1991_buf_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(58)); -- 
    -- CP-element group 59:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_sample_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_sample_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_update_start__ps
      -- CP-element group 60: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_3269_elements(61) <= nicRxFromMacDaemon_CP_3269_elements(62);
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	61 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/type_cast_1993_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_3269_elements(60), ack => nicRxFromMacDaemon_CP_3269_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	25 
    -- CP-element group 63: 	43 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_start/req
      -- CP-element group 63: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_sample_start_
      -- 
    req_3521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(63), ack => MUX_2021_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(25) & nicRxFromMacDaemon_CP_3269_elements(43) & nicRxFromMacDaemon_CP_3269_elements(65);
      gj_nicRxFromMacDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	68 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_complete/req
      -- 
    req_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(64), ack => MUX_2021_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(66) & nicRxFromMacDaemon_CP_3269_elements(68);
      gj_nicRxFromMacDaemon_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	23 
    -- CP-element group 65: 	39 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_start/ack
      -- CP-element group 65: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_sample_completed_
      -- 
    ack_3522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2021_inst_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/MUX_2021_complete/ack
      -- 
    ack_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_2021_inst_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	66 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Sample/$entry
      -- 
    req_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(67), ack => WPIPE_nic_rx_to_header_2012_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(25) & nicRxFromMacDaemon_CP_3269_elements(66) & nicRxFromMacDaemon_CP_3269_elements(69);
      gj_nicRxFromMacDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	23 
    -- CP-element group 68: 	64 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Update/req
      -- 
    ack_3536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_2012_inst_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(68)); -- 
    req_3540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(68), ack => WPIPE_nic_rx_to_header_2012_inst_req_1); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	78 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Update/ack
      -- CP-element group 69: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_header_2012_Update/$exit
      -- 
    ack_3541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_2012_inst_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	43 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Sample/req
      -- CP-element group 70: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Sample/$entry
      -- 
    req_3549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(70), ack => WPIPE_nic_rx_to_packet_2023_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(43) & nicRxFromMacDaemon_CP_3269_elements(72);
      gj_nicRxFromMacDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	39 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Update/req
      -- CP-element group 71: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Sample/$exit
      -- 
    ack_3550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_2023_inst_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(71)); -- 
    req_3554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(71), ack => WPIPE_nic_rx_to_packet_2023_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	78 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/WPIPE_nic_rx_to_packet_2023_update_completed_
      -- 
    ack_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_2023_inst_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	25 
    -- CP-element group 73: 	43 
    -- CP-element group 73: 	49 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Sample/crr
      -- CP-element group 73: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_sample_start_
      -- 
    crr_3563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(73), ack => call_stmt_2049_call_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(25) & nicRxFromMacDaemon_CP_3269_elements(43) & nicRxFromMacDaemon_CP_3269_elements(49) & nicRxFromMacDaemon_CP_3269_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Update/ccr
      -- 
    ccr_3568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(74), ack => call_stmt_2049_call_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicRxFromMacDaemon_CP_3269_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	23 
    -- CP-element group 75: 	39 
    -- CP-element group 75: 	45 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Sample/cra
      -- CP-element group 75: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_sample_completed_
      -- 
    cra_3564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2049_call_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/call_stmt_2049_Update/cca
      -- 
    cca_3569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2049_call_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(76)); -- 
    -- CP-element group 77:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	16 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	17 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_3269_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_3269_elements(16), ack => nicRxFromMacDaemon_CP_3269_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	19 
    -- CP-element group 78: 	69 
    -- CP-element group 78: 	72 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	13 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1949/do_while_stmt_1980/do_while_stmt_1980_loop_body/$exit
      -- 
    nicRxFromMacDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_3269_elements(19) & nicRxFromMacDaemon_CP_3269_elements(69) & nicRxFromMacDaemon_CP_3269_elements(72) & nicRxFromMacDaemon_CP_3269_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	12 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_exit/$exit
      -- CP-element group 79: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_exit/ack
      -- 
    ack_3574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1980_branch_ack_0, ack => nicRxFromMacDaemon_CP_3269_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	12 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_taken/$exit
      -- CP-element group 80: 	 branch_block_stmt_1949/do_while_stmt_1980/loop_taken/ack
      -- 
    ack_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1980_branch_ack_1, ack => nicRxFromMacDaemon_CP_3269_elements(80)); -- 
    -- CP-element group 81:  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	10 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	2 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1949/do_while_stmt_1980/$exit
      -- 
    nicRxFromMacDaemon_CP_3269_elements(81) <= nicRxFromMacDaemon_CP_3269_elements(10);
    -- CP-element group 82:  merge  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	0 
    -- CP-element group 82: 	2 
    -- CP-element group 82: 	5 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	3 
    -- CP-element group 82: 	4 
    -- CP-element group 82:  members (13) 
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/$entry
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961__entry__
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Update/ccr
      -- CP-element group 82: 	 branch_block_stmt_1949/merge_stmt_1951__exit__
      -- CP-element group 82: 	 branch_block_stmt_1949/merge_stmt_1951_PhiAck/$entry
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Sample/crr
      -- CP-element group 82: 	 branch_block_stmt_1949/call_stmt_1961/call_stmt_1961_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1949/merge_stmt_1951_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_1949/merge_stmt_1951_PhiAck/dummy
      -- CP-element group 82: 	 branch_block_stmt_1949/merge_stmt_1951_PhiAck/$exit
      -- 
    ccr_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(82), ack => call_stmt_1961_call_req_1); -- 
    crr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_3269_elements(82), ack => call_stmt_1961_call_req_0); -- 
    nicRxFromMacDaemon_CP_3269_elements(82) <= OrReduce(nicRxFromMacDaemon_CP_3269_elements(0) & nicRxFromMacDaemon_CP_3269_elements(2) & nicRxFromMacDaemon_CP_3269_elements(5));
    nicRxFromMacDaemon_do_while_stmt_1980_terminator_3579: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_1980_terminator_3579", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_3269_elements(13),loop_continue => nicRxFromMacDaemon_CP_3269_elements(80),loop_terminate => nicRxFromMacDaemon_CP_3269_elements(79),loop_back => nicRxFromMacDaemon_CP_3269_elements(11),loop_exit => nicRxFromMacDaemon_CP_3269_elements(10),clk => clk, reset => reset); -- 
    phi_stmt_1982_phi_seq_3451_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_3269_elements(26);
      nicRxFromMacDaemon_CP_3269_elements(31)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_3269_elements(33);
      nicRxFromMacDaemon_CP_3269_elements(32)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_3269_elements(34);
      nicRxFromMacDaemon_CP_3269_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_3269_elements(28);
      nicRxFromMacDaemon_CP_3269_elements(35)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_3269_elements(35);
      nicRxFromMacDaemon_CP_3269_elements(36)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_3269_elements(37);
      nicRxFromMacDaemon_CP_3269_elements(29) <= phi_mux_reqs(1);
      phi_stmt_1982_phi_seq_3451 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1982_phi_seq_3451") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_3269_elements(18), 
          phi_sample_ack => nicRxFromMacDaemon_CP_3269_elements(24), 
          phi_update_req => nicRxFromMacDaemon_CP_3269_elements(20), 
          phi_update_ack => nicRxFromMacDaemon_CP_3269_elements(25), 
          phi_mux_ack => nicRxFromMacDaemon_CP_3269_elements(30), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1989_phi_seq_3513_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_3269_elements(50);
      nicRxFromMacDaemon_CP_3269_elements(55)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_3269_elements(57);
      nicRxFromMacDaemon_CP_3269_elements(56)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_3269_elements(58);
      nicRxFromMacDaemon_CP_3269_elements(51) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_3269_elements(52);
      nicRxFromMacDaemon_CP_3269_elements(59)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_3269_elements(59);
      nicRxFromMacDaemon_CP_3269_elements(60)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_3269_elements(61);
      nicRxFromMacDaemon_CP_3269_elements(53) <= phi_mux_reqs(1);
      phi_stmt_1989_phi_seq_3513 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1989_phi_seq_3513") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_3269_elements(46), 
          phi_sample_ack => nicRxFromMacDaemon_CP_3269_elements(47), 
          phi_update_req => nicRxFromMacDaemon_CP_3269_elements(48), 
          phi_update_ack => nicRxFromMacDaemon_CP_3269_elements(49), 
          phi_mux_ack => nicRxFromMacDaemon_CP_3269_elements(54), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3403_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_3269_elements(14);
        preds(1)  <= nicRxFromMacDaemon_CP_3269_elements(15);
        entry_tmerge_3403 : transition_merge -- 
          generic map(name => " entry_tmerge_3403")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_3269_elements(16));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_2036_wire : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_1965_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2056_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u65_u73_2019_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_2005_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2008_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2015_wire : std_logic_vector(0 downto 0);
    signal LSTATE_1982 : std_logic_vector(1 downto 0);
    signal MUX_2021_wire : std_logic_vector(72 downto 0);
    signal NOT_u1_u1_1966_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1956_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1974_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_2045_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1963_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_2054_wire : std_logic_vector(31 downto 0);
    signal RPIPE_mac_to_nic_data_1988_wire : std_logic_vector(72 downto 0);
    signal RX_1986 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_2018_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_1985_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_2004_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_2028_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_2007_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_2014_wire_constant : std_logic_vector(1 downto 0);
    signal ignore_resp0_1961 : std_logic_vector(31 downto 0);
    signal ignore_resp1_1979 : std_logic_vector(31 downto 0);
    signal ignore_resp2_2049 : std_logic_vector(31 downto 0);
    signal konst_1957_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1964_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1975_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2046_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2055_wire_constant : std_logic_vector(31 downto 0);
    signal nLSTATE_2001 : std_logic_vector(1 downto 0);
    signal nLSTATE_2001_1984_buffered : std_logic_vector(1 downto 0);
    signal npkt_cnt_2039 : std_logic_vector(31 downto 0);
    signal npkt_cnt_2039_1991_buffered : std_logic_vector(31 downto 0);
    signal pkt_cnt_1989 : std_logic_vector(31 downto 0);
    signal pkt_complete_2030 : std_logic_vector(0 downto 0);
    signal slice_2017_wire : std_logic_vector(64 downto 0);
    signal type_cast_1953_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1959_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1971_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1977_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1993_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2035_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2042_wire_constant : std_logic_vector(0 downto 0);
    signal write_to_header_2010 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1956_wire_constant <= "1111";
    NOT_u4_u4_1974_wire_constant <= "1111";
    NOT_u4_u4_2045_wire_constant <= "1111";
    R_HEADER_TKEEP_2018_wire_constant <= "00111111";
    R_S0_1985_wire_constant <= "00";
    R_S0_2004_wire_constant <= "00";
    R_S0_2028_wire_constant <= "00";
    R_S1_2007_wire_constant <= "01";
    R_S1_2014_wire_constant <= "01";
    konst_1957_wire_constant <= "010110";
    konst_1964_wire_constant <= "00000000000000000000000000000000";
    konst_1975_wire_constant <= "010110";
    konst_2046_wire_constant <= "010111";
    konst_2055_wire_constant <= "00000000000000000000000000000000";
    type_cast_1953_wire_constant <= "0";
    type_cast_1959_wire_constant <= "00000000000000000000000000000000";
    type_cast_1971_wire_constant <= "0";
    type_cast_1977_wire_constant <= "00000000000000000000000000000001";
    type_cast_1993_wire_constant <= "00000000000000000000000000000000";
    type_cast_2035_wire_constant <= "00000000000000000000000000000001";
    type_cast_2042_wire_constant <= "0";
    phi_stmt_1982: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nLSTATE_2001_1984_buffered & R_S0_1985_wire_constant;
      req <= phi_stmt_1982_req_0 & phi_stmt_1982_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1982",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1982_ack_0,
          idata => idata,
          odata => LSTATE_1982,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1982
    phi_stmt_1989: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= npkt_cnt_2039_1991_buffered & type_cast_1993_wire_constant;
      req <= phi_stmt_1989_req_0 & phi_stmt_1989_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1989",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1989_ack_0,
          idata => idata,
          odata => pkt_cnt_1989,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1989
    MUX_2021_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_2021_inst_req_0;
      MUX_2021_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_2021_inst_req_1;
      MUX_2021_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_2010(0);
      MUX_2021_inst_gI: SplitGuardInterface generic map(name => "MUX_2021_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_2021_inst: SelectSplitProtocol generic map(name => "MUX_2021_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_2019_wire, y => RX_1986, sel => EQ_u2_u1_2015_wire, z => MUX_2021_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_2038_inst
    npkt_cnt_2039 <= ADD_u32_u32_2036_wire when (pkt_complete_2030(0) /=  '0') else pkt_cnt_1989;
    -- flow-through slice operator slice_2017_inst
    slice_2017_wire <= RX_1986(72 downto 8);
    nLSTATE_2001_1984_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_2001_1984_buf_req_0;
      nLSTATE_2001_1984_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_2001_1984_buf_req_1;
      nLSTATE_2001_1984_buf_ack_1<= rack(0);
      nLSTATE_2001_1984_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_2001_1984_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_2001,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_2001_1984_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_2039_1991_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_2039_1991_buf_req_0;
      npkt_cnt_2039_1991_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_2039_1991_buf_req_1;
      npkt_cnt_2039_1991_buf_ack_1<= rack(0);
      npkt_cnt_2039_1991_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_2039_1991_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_2039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_2039_1991_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1986
    process(RPIPE_mac_to_nic_data_1988_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_1988_wire(72 downto 0);
      RX_1986 <= tmp_var; -- 
    end process;
    do_while_stmt_1980_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_2056_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1980_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1980_branch_req_0,
          ack0 => do_while_stmt_1980_branch_ack_0,
          ack1 => do_while_stmt_1980_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1962_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1966_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1962_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1962_branch_req_0,
          ack0 => if_stmt_1962_branch_ack_0,
          ack1 => if_stmt_1962_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_2036_inst
    process(pkt_cnt_1989) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pkt_cnt_1989, type_cast_2035_wire_constant, tmp_var);
      ADD_u32_u32_2036_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1965_inst
    process(RPIPE_CONTROL_REGISTER_1963_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1963_wire, konst_1964_wire_constant, tmp_var);
      BITSEL_u32_u1_1965_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_2056_inst
    process(RPIPE_CONTROL_REGISTER_2054_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_2054_wire, konst_2055_wire_constant, tmp_var);
      BITSEL_u32_u1_2056_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u65_u73_2019_inst
    process(slice_2017_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_2017_wire, R_HEADER_TKEEP_2018_wire_constant, tmp_var);
      CONCAT_u65_u73_2019_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2005_inst
    process(LSTATE_1982) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1982, R_S0_2004_wire_constant, tmp_var);
      EQ_u2_u1_2005_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2008_inst
    process(LSTATE_1982) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1982, R_S1_2007_wire_constant, tmp_var);
      EQ_u2_u1_2008_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2015_inst
    process(LSTATE_1982) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1982, R_S1_2014_wire_constant, tmp_var);
      EQ_u2_u1_2015_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2029_inst
    process(nLSTATE_2001) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(nLSTATE_2001, R_S0_2028_wire_constant, tmp_var);
      pkt_complete_2030 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1966_inst
    process(BITSEL_u32_u1_1965_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1965_wire, tmp_var);
      NOT_u1_u1_1966_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2009_inst
    process(EQ_u2_u1_2005_wire, EQ_u2_u1_2008_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_2005_wire, EQ_u2_u1_2008_wire, tmp_var);
      write_to_header_2010 <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1963_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_2054_wire <= CONTROL_REGISTER;
    -- shared inport operator group (2) : RPIPE_mac_to_nic_data_1988_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_1988_inst_req_0;
      RPIPE_mac_to_nic_data_1988_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_1988_inst_req_1;
      RPIPE_mac_to_nic_data_1988_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_1988_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_2_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_2: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_2", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_2012_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_2012_inst_req_0;
      WPIPE_nic_rx_to_header_2012_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_2012_inst_req_1;
      WPIPE_nic_rx_to_header_2012_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_2010(0);
      data_in <= MUX_2021_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_2023_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_2023_inst_req_0;
      WPIPE_nic_rx_to_packet_2023_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_2023_inst_req_1;
      WPIPE_nic_rx_to_packet_2023_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_1986;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1961_call call_stmt_1979_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1961_call_req_0;
      reqL_unguarded(0) <= call_stmt_1979_call_req_0;
      call_stmt_1961_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1979_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1961_call_req_1;
      reqR_unguarded(0) <= call_stmt_1979_call_req_1;
      call_stmt_1961_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1979_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      AccessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1953_wire_constant & NOT_u4_u4_1956_wire_constant & konst_1957_wire_constant & type_cast_1959_wire_constant & type_cast_1971_wire_constant & NOT_u4_u4_1974_wire_constant & konst_1975_wire_constant & type_cast_1977_wire_constant;
      ignore_resp0_1961 <= data_out(63 downto 32);
      ignore_resp1_1979 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(1),
          ackR => AccessRegister_call_acks(1),
          dataR => AccessRegister_call_data(85 downto 43),
          tagR => AccessRegister_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(1), -- cross-over
          ackL => AccessRegister_return_reqs(1), -- cross-over
          dataL => AccessRegister_return_data(63 downto 32),
          tagL => AccessRegister_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_nextLSTATE_5243: nextLSTATE_Volatile port map(RX => RX_1986, LSTATE => LSTATE_1982, nLSTATE => nLSTATE_2001); 
    -- shared call operator group (2) : call_stmt_2049_call 
    AccessRegister_call_group_2: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2049_call_req_0;
      call_stmt_2049_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2049_call_req_1;
      call_stmt_2049_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= pkt_complete_2030(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_2_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2042_wire_constant & NOT_u4_u4_2045_wire_constant & konst_2046_wire_constant & pkt_cnt_1989;
      ignore_resp2_2049 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(35 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(67 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(31 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(35 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
    updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(35 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 37)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_944_start: Boolean;
  signal popFromQueue_CP_944_symbol: Boolean;
  -- volatile/operator module components. 
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_955_call_req_0 : boolean;
  signal call_stmt_955_call_ack_0 : boolean;
  signal call_stmt_955_call_req_1 : boolean;
  signal call_stmt_955_call_ack_1 : boolean;
  signal call_stmt_969_call_req_0 : boolean;
  signal call_stmt_969_call_ack_0 : boolean;
  signal call_stmt_969_call_req_1 : boolean;
  signal call_stmt_969_call_ack_1 : boolean;
  signal call_stmt_974_call_req_0 : boolean;
  signal call_stmt_974_call_ack_0 : boolean;
  signal call_stmt_974_call_req_1 : boolean;
  signal call_stmt_974_call_ack_1 : boolean;
  signal call_stmt_982_call_req_0 : boolean;
  signal call_stmt_982_call_ack_0 : boolean;
  signal call_stmt_982_call_req_1 : boolean;
  signal call_stmt_982_call_ack_1 : boolean;
  signal call_stmt_985_call_req_0 : boolean;
  signal call_stmt_985_call_ack_0 : boolean;
  signal call_stmt_985_call_req_1 : boolean;
  signal call_stmt_985_call_ack_1 : boolean;
  signal call_stmt_1005_call_req_0 : boolean;
  signal call_stmt_1005_call_ack_0 : boolean;
  signal call_stmt_1005_call_req_1 : boolean;
  signal call_stmt_1005_call_ack_1 : boolean;
  signal call_stmt_1010_call_req_0 : boolean;
  signal call_stmt_1010_call_ack_0 : boolean;
  signal call_stmt_1010_call_req_1 : boolean;
  signal call_stmt_1010_call_ack_1 : boolean;
  signal call_stmt_1017_call_req_0 : boolean;
  signal call_stmt_1017_call_ack_0 : boolean;
  signal call_stmt_1017_call_req_1 : boolean;
  signal call_stmt_1017_call_ack_1 : boolean;
  signal call_stmt_1028_call_req_0 : boolean;
  signal call_stmt_1028_call_ack_0 : boolean;
  signal call_stmt_1028_call_req_1 : boolean;
  signal call_stmt_1028_call_ack_1 : boolean;
  signal W_status_1029_inst_req_0 : boolean;
  signal W_status_1029_inst_ack_0 : boolean;
  signal W_status_1029_inst_req_1 : boolean;
  signal W_status_1029_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 37) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(tag_length + 36 downto 37) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 36 downto 37);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_944_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_944_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_944_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_944_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_944: Block -- control-path 
    signal popFromQueue_CP_944_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_944_elements(0) <= popFromQueue_CP_944_start;
    popFromQueue_CP_944_symbol <= popFromQueue_CP_944_elements(24);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/$entry
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_sample_start_
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_update_start_
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Sample/$entry
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Sample/crr
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Update/$entry
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Update/ccr
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_update_start_
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Update/$entry
      -- CP-element group 0: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Update/ccr
      -- 
    crr_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(0), ack => call_stmt_955_call_req_0); -- 
    ccr_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(0), ack => call_stmt_955_call_req_1); -- 
    ccr_976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(0), ack => call_stmt_969_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_sample_completed_
      -- CP-element group 1: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Sample/$exit
      -- CP-element group 1: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Sample/cra
      -- 
    cra_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_955_call_ack_0, ack => popFromQueue_CP_944_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_update_completed_
      -- CP-element group 2: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Update/$exit
      -- CP-element group 2: 	 call_stmt_955_to_call_stmt_969/call_stmt_955_Update/cca
      -- CP-element group 2: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_sample_start_
      -- CP-element group 2: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Sample/$entry
      -- CP-element group 2: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Sample/crr
      -- 
    cca_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_955_call_ack_1, ack => popFromQueue_CP_944_elements(2)); -- 
    crr_971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(2), ack => call_stmt_969_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_sample_completed_
      -- CP-element group 3: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Sample/$exit
      -- CP-element group 3: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Sample/cra
      -- 
    cra_972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_969_call_ack_0, ack => popFromQueue_CP_944_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	13 
    -- CP-element group 4: 	16 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (26) 
      -- CP-element group 4: 	 call_stmt_955_to_call_stmt_969/$exit
      -- CP-element group 4: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_update_completed_
      -- CP-element group 4: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Update/$exit
      -- CP-element group 4: 	 call_stmt_955_to_call_stmt_969/call_stmt_969_Update/cca
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_sample_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_update_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Sample/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Sample/crr
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Update/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Update/ccr
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_update_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Update/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Update/ccr
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_update_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Update/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Update/ccr
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_update_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Update/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Update/ccr
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_update_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Update/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Update/ccr
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_update_start_
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Update/$entry
      -- CP-element group 4: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Update/ccr
      -- 
    cca_977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_969_call_ack_1, ack => popFromQueue_CP_944_elements(4)); -- 
    crr_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_974_call_req_0); -- 
    ccr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_974_call_req_1); -- 
    ccr_1007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_982_call_req_1); -- 
    ccr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_985_call_req_1); -- 
    ccr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_1005_call_req_1); -- 
    ccr_1049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_1010_call_req_1); -- 
    ccr_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(4), ack => call_stmt_1017_call_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_sample_completed_
      -- CP-element group 5: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Sample/$exit
      -- CP-element group 5: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Sample/cra
      -- 
    cra_989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_974_call_ack_0, ack => popFromQueue_CP_944_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	11 
    -- CP-element group 6: 	14 
    -- CP-element group 6: 	17 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_update_completed_
      -- CP-element group 6: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Update/$exit
      -- CP-element group 6: 	 call_stmt_974_to_call_stmt_1017/call_stmt_974_Update/cca
      -- CP-element group 6: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_sample_start_
      -- CP-element group 6: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Sample/$entry
      -- CP-element group 6: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Sample/crr
      -- 
    cca_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_974_call_ack_1, ack => popFromQueue_CP_944_elements(6)); -- 
    crr_1002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(6), ack => call_stmt_982_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_sample_completed_
      -- CP-element group 7: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Sample/$exit
      -- CP-element group 7: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Sample/cra
      -- 
    cra_1003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_982_call_ack_0, ack => popFromQueue_CP_944_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_update_completed_
      -- CP-element group 8: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Update/$exit
      -- CP-element group 8: 	 call_stmt_974_to_call_stmt_1017/call_stmt_982_Update/cca
      -- CP-element group 8: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_sample_start_
      -- CP-element group 8: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Sample/$entry
      -- CP-element group 8: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Sample/crr
      -- 
    cca_1008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_982_call_ack_1, ack => popFromQueue_CP_944_elements(8)); -- 
    crr_1016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(8), ack => call_stmt_985_call_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_sample_completed_
      -- CP-element group 9: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Sample/$exit
      -- CP-element group 9: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Sample/cra
      -- 
    cra_1017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_985_call_ack_0, ack => popFromQueue_CP_944_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	17 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_update_completed_
      -- CP-element group 10: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Update/$exit
      -- CP-element group 10: 	 call_stmt_974_to_call_stmt_1017/call_stmt_985_Update/cca
      -- 
    cca_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_985_call_ack_1, ack => popFromQueue_CP_944_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_sample_start_
      -- CP-element group 11: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Sample/$entry
      -- CP-element group 11: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Sample/crr
      -- 
    crr_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(11), ack => call_stmt_1005_call_req_0); -- 
    popFromQueue_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_944_elements(6) & popFromQueue_CP_944_elements(10);
      gj_popFromQueue_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_944_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_sample_completed_
      -- CP-element group 12: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Sample/$exit
      -- CP-element group 12: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Sample/cra
      -- 
    cra_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1005_call_ack_0, ack => popFromQueue_CP_944_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	4 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_update_completed_
      -- CP-element group 13: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Update/$exit
      -- CP-element group 13: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1005_Update/cca
      -- 
    cca_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1005_call_ack_1, ack => popFromQueue_CP_944_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: 	8 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_sample_start_
      -- CP-element group 14: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Sample/$entry
      -- CP-element group 14: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Sample/crr
      -- 
    crr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(14), ack => call_stmt_1010_call_req_0); -- 
    popFromQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= popFromQueue_CP_944_elements(6) & popFromQueue_CP_944_elements(8) & popFromQueue_CP_944_elements(13);
      gj_popFromQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_944_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_sample_completed_
      -- CP-element group 15: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Sample/$exit
      -- CP-element group 15: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Sample/cra
      -- 
    cra_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1010_call_ack_0, ack => popFromQueue_CP_944_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	4 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_update_completed_
      -- CP-element group 16: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Update/$exit
      -- CP-element group 16: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1010_Update/cca
      -- 
    cca_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1010_call_ack_1, ack => popFromQueue_CP_944_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	6 
    -- CP-element group 17: 	10 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_sample_start_
      -- CP-element group 17: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Sample/$entry
      -- CP-element group 17: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Sample/crr
      -- 
    crr_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(17), ack => call_stmt_1017_call_req_0); -- 
    popFromQueue_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= popFromQueue_CP_944_elements(6) & popFromQueue_CP_944_elements(10) & popFromQueue_CP_944_elements(16);
      gj_popFromQueue_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_944_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_sample_completed_
      -- CP-element group 18: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Sample/$exit
      -- CP-element group 18: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Sample/cra
      -- 
    cra_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1017_call_ack_0, ack => popFromQueue_CP_944_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (17) 
      -- CP-element group 19: 	 call_stmt_974_to_call_stmt_1017/$exit
      -- CP-element group 19: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_update_completed_
      -- CP-element group 19: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Update/$exit
      -- CP-element group 19: 	 call_stmt_974_to_call_stmt_1017/call_stmt_1017_Update/cca
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/$entry
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_sample_start_
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_update_start_
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Sample/crr
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Update/$entry
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Update/ccr
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_sample_start_
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_update_start_
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Sample/req
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Update/$entry
      -- CP-element group 19: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Update/req
      -- 
    cca_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1017_call_ack_1, ack => popFromQueue_CP_944_elements(19)); -- 
    crr_1075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(19), ack => call_stmt_1028_call_req_0); -- 
    ccr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(19), ack => call_stmt_1028_call_req_1); -- 
    req_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(19), ack => W_status_1029_inst_req_0); -- 
    req_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_944_elements(19), ack => W_status_1029_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_sample_completed_
      -- CP-element group 20: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Sample/cra
      -- 
    cra_1076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1028_call_ack_0, ack => popFromQueue_CP_944_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_update_completed_
      -- CP-element group 21: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Update/$exit
      -- CP-element group 21: 	 call_stmt_1028_to_assign_stmt_1031/call_stmt_1028_Update/cca
      -- 
    cca_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1028_call_ack_1, ack => popFromQueue_CP_944_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_sample_completed_
      -- CP-element group 22: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Sample/$exit
      -- CP-element group 22: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Sample/ack
      -- 
    ack_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1029_inst_ack_0, ack => popFromQueue_CP_944_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_update_completed_
      -- CP-element group 23: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Update/$exit
      -- CP-element group 23: 	 call_stmt_1028_to_assign_stmt_1031/assign_stmt_1031_Update/ack
      -- 
    ack_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1029_inst_ack_1, ack => popFromQueue_CP_944_elements(23)); -- 
    -- CP-element group 24:  join  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 $exit
      -- CP-element group 24: 	 call_stmt_1028_to_assign_stmt_1031/$exit
      -- 
    popFromQueue_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_944_elements(23) & popFromQueue_CP_944_elements(21);
      gj_popFromQueue_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_944_elements(24), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_998_wire : std_logic_vector(31 downto 0);
    signal ADD_u36_u36_951_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_948_wire_constant : std_logic_vector(7 downto 0);
    signal Queue_Length_982 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1016_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_990_wire : std_logic_vector(31 downto 0);
    signal ba_and_misc_955 : std_logic_vector(63 downto 0);
    signal konst_950_wire_constant : std_logic_vector(35 downto 0);
    signal konst_989_wire_constant : std_logic_vector(31 downto 0);
    signal konst_995_wire_constant : std_logic_vector(31 downto 0);
    signal konst_997_wire_constant : std_logic_vector(31 downto 0);
    signal lock_n_965 : std_logic_vector(0 downto 0);
    signal m_ok_969 : std_logic_vector(0 downto 0);
    signal misc_959 : std_logic_vector(31 downto 0);
    signal next_ri_1000 : std_logic_vector(31 downto 0);
    signal q_empty_979 : std_logic_vector(0 downto 0);
    signal read_index_974 : std_logic_vector(31 downto 0);
    signal round_off_992 : std_logic_vector(0 downto 0);
    signal total_msgs_985 : std_logic_vector(31 downto 0);
    signal type_cast_1015_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_945_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_953_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_963_wire_constant : std_logic_vector(31 downto 0);
    signal write_index_974 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_948_wire_constant <= "11111111";
    konst_950_wire_constant <= "000000000000000000000000000000011000";
    konst_989_wire_constant <= "00000000000000000000000000000001";
    konst_995_wire_constant <= "00000000000000000000000000000000";
    konst_997_wire_constant <= "00000000000000000000000000000001";
    type_cast_1015_wire_constant <= "00000000000000000000000000000001";
    type_cast_943_wire_constant <= "0";
    type_cast_945_wire_constant <= "1";
    type_cast_953_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_963_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_999_inst
    next_ri_1000 <= konst_995_wire_constant when (round_off_992(0) /=  '0') else ADD_u32_u32_998_wire;
    -- flow-through slice operator slice_958_inst
    misc_959 <= ba_and_misc_955(31 downto 0);
    W_status_1029_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_1029_inst_req_0;
      W_status_1029_inst_ack_0<= wack(0);
      rreq(0) <= W_status_1029_inst_req_1;
      W_status_1029_inst_ack_1<= rack(0);
      W_status_1029_inst : InterlockBuffer generic map ( -- 
        name => "W_status_1029_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_empty_979,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator ADD_u32_u32_998_inst
    process(read_index_974) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_index_974, konst_997_wire_constant, tmp_var);
      ADD_u32_u32_998_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_951_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_950_wire_constant, tmp_var);
      ADD_u36_u36_951_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_964_inst
    process(misc_959) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(misc_959, type_cast_963_wire_constant, tmp_var);
      lock_n_965 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_978_inst
    process(write_index_974, read_index_974) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_974, read_index_974, tmp_var);
      q_empty_979 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_991_inst
    process(read_index_974, SUB_u32_u32_990_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(read_index_974, SUB_u32_u32_990_wire, tmp_var);
      round_off_992 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1016_inst
    process(total_msgs_985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(total_msgs_985, type_cast_1015_wire_constant, tmp_var);
      SUB_u32_u32_1016_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_990_inst
    process(Queue_Length_982) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(Queue_Length_982, konst_989_wire_constant, tmp_var);
      SUB_u32_u32_990_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1005_call 
    getQueueElement_call_group_0: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1005_call_req_0;
      call_stmt_1005_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1005_call_req_1;
      call_stmt_1005_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_979(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_0_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & read_index_974;
      q_r_data_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(67 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(31 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1010_call 
    setQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1010_call_req_0;
      call_stmt_1010_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1010_call_req_1;
      call_stmt_1010_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_979(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_index_974 & next_ri_1000;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1017_call 
    updateTotalMessages_call_group_2: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1017_call_req_0;
      call_stmt_1017_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1017_call_req_1;
      call_stmt_1017_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_979(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateTotalMessages_call_group_2_gI: SplitGuardInterface generic map(name => "updateTotalMessages_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & SUB_u32_u32_1016_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateTotalMessages_call_reqs(0),
          ackR => updateTotalMessages_call_acks(0),
          dataR => updateTotalMessages_call_data(67 downto 0),
          tagR => updateTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => updateTotalMessages_return_acks(0), -- cross-over
          ackL => updateTotalMessages_return_reqs(0), -- cross-over
          tagL => updateTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1028_call 
    releaseLock_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1028_call_req_0;
      call_stmt_1028_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1028_call_req_1;
      call_stmt_1028_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_965(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_3_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(35 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_955_call 
    accessMemory_call_group_4: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_955_call_req_0;
      call_stmt_955_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_955_call_req_1;
      call_stmt_955_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_4_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_943_wire_constant & type_cast_945_wire_constant & NOT_u8_u8_948_wire_constant & ADD_u36_u36_951_wire & type_cast_953_wire_constant;
      ba_and_misc_955 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_969_call 
    acquireLock_call_group_5: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_969_call_req_0;
      call_stmt_969_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_969_call_req_1;
      call_stmt_969_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_965(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_5_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_969 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(35 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_974_call 
    getQueuePointers_call_group_6: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_974_call_req_0;
      call_stmt_974_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_974_call_req_1;
      call_stmt_974_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_6_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_index_974 <= data_out(63 downto 32);
      read_index_974 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_982_call 
    getQueueLength_call_group_7: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_982_call_req_0;
      call_stmt_982_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_982_call_req_1;
      call_stmt_982_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_7_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      Queue_Length_982 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(35 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_985_call 
    getTotalMessages_call_group_8: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_985_call_req_0;
      call_stmt_985_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_985_call_req_1;
      call_stmt_985_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_8_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      total_msgs_985 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(35 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_1799_start: Boolean;
  signal populateRxQueue_CP_1799_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(31 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1448_call_req_0 : boolean;
  signal call_stmt_1448_call_ack_0 : boolean;
  signal call_stmt_1448_call_req_1 : boolean;
  signal call_stmt_1448_call_ack_1 : boolean;
  signal call_stmt_1465_call_req_0 : boolean;
  signal call_stmt_1465_call_ack_0 : boolean;
  signal call_stmt_1465_call_req_1 : boolean;
  signal call_stmt_1465_call_ack_1 : boolean;
  signal AND_u6_u6_1474_inst_req_0 : boolean;
  signal AND_u6_u6_1474_inst_ack_0 : boolean;
  signal AND_u6_u6_1474_inst_req_1 : boolean;
  signal AND_u6_u6_1474_inst_ack_1 : boolean;
  signal if_stmt_1479_branch_req_0 : boolean;
  signal if_stmt_1479_branch_ack_1 : boolean;
  signal if_stmt_1479_branch_ack_0 : boolean;
  signal call_stmt_1484_call_req_0 : boolean;
  signal call_stmt_1484_call_ack_0 : boolean;
  signal call_stmt_1484_call_req_1 : boolean;
  signal call_stmt_1484_call_ack_1 : boolean;
  signal if_stmt_1485_branch_req_0 : boolean;
  signal if_stmt_1485_branch_ack_1 : boolean;
  signal if_stmt_1485_branch_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_ack_1 : boolean;
  signal AND_u6_u6_1426_inst_req_0 : boolean;
  signal AND_u6_u6_1426_inst_ack_0 : boolean;
  signal AND_u6_u6_1426_inst_req_1 : boolean;
  signal AND_u6_u6_1426_inst_ack_1 : boolean;
  signal phi_stmt_1417_req_0 : boolean;
  signal n_q_index_1475_1427_buf_req_0 : boolean;
  signal n_q_index_1475_1427_buf_ack_0 : boolean;
  signal n_q_index_1475_1427_buf_req_1 : boolean;
  signal n_q_index_1475_1427_buf_ack_1 : boolean;
  signal phi_stmt_1417_req_1 : boolean;
  signal phi_stmt_1417_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_1799_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1799_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_1799_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1799_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_1799: Block -- control-path 
    signal populateRxQueue_CP_1799_elements: BooleanArray(25 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_1799_elements(0) <= populateRxQueue_CP_1799_start;
    populateRxQueue_CP_1799_symbol <= populateRxQueue_CP_1799_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1415/$entry
      -- CP-element group 0: 	 branch_block_stmt_1415/branch_block_stmt_1415__entry__
      -- CP-element group 0: 	 branch_block_stmt_1415/merge_stmt_1416__entry__
      -- CP-element group 0: 	 branch_block_stmt_1415/merge_stmt_1416_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1415/$exit
      -- CP-element group 1: 	 branch_block_stmt_1415/branch_block_stmt_1415__exit__
      -- CP-element group 1: 	 branch_block_stmt_1415/if_stmt_1479__exit__
      -- 
    populateRxQueue_CP_1799_elements(1) <= OrReduce(populateRxQueue_CP_1799_elements(14) & populateRxQueue_CP_1799_elements(16));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	25 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Sample/cra
      -- 
    cra_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1448_call_ack_0, ack => populateRxQueue_CP_1799_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	25 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Sample/crr
      -- 
    cca_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1448_call_ack_1, ack => populateRxQueue_CP_1799_elements(3)); -- 
    crr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(3), ack => call_stmt_1465_call_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Sample/cra
      -- 
    cra_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1465_call_ack_0, ack => populateRxQueue_CP_1799_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Update/cca
      -- 
    cca_1843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1465_call_ack_1, ack => populateRxQueue_CP_1799_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	25 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Sample/ra
      -- 
    ra_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1474_inst_ack_0, ack => populateRxQueue_CP_1799_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	25 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Update/ca
      -- 
    ca_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1474_inst_ack_1, ack => populateRxQueue_CP_1799_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (22) 
      -- CP-element group 8: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475__exit__
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479__entry__
      -- CP-element group 8: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/$exit
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/$exit
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/NOT_u1_u1_1481/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_1415/NOT_u1_u1_1481_place
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_1415/if_stmt_1479_else_link/$entry
      -- 
    branch_req_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(8), ack => if_stmt_1479_branch_req_0); -- 
    populateRxQueue_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "populateRxQueue_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1799_elements(5) & populateRxQueue_CP_1799_elements(7);
      gj_populateRxQueue_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1799_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_1415/if_stmt_1479_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_1415/if_stmt_1479_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484__entry__
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/$entry
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Update/ccr
      -- 
    if_choice_transition_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1479_branch_ack_1, ack => populateRxQueue_CP_1799_elements(9)); -- 
    crr_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(9), ack => call_stmt_1484_call_req_0); -- 
    ccr_1910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(9), ack => call_stmt_1484_call_req_1); -- 
    -- CP-element group 10:  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_1415/if_stmt_1479_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_1415/if_stmt_1479_else_link/else_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_1415/assign_stmt_1494__entry__
      -- CP-element group 10: 	 branch_block_stmt_1415/assign_stmt_1494/$entry
      -- CP-element group 10: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Sample/req
      -- 
    else_choice_transition_1890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1479_branch_ack_0, ack => populateRxQueue_CP_1799_elements(10)); -- 
    req_1961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(10), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Sample/cra
      -- 
    cra_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1484_call_ack_0, ack => populateRxQueue_CP_1799_elements(11)); -- 
    -- CP-element group 12:  branch  transition  place  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (27) 
      -- CP-element group 12: 	 branch_block_stmt_1415/call_stmt_1484__exit__
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485__entry__
      -- CP-element group 12: 	 branch_block_stmt_1415/call_stmt_1484/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/call_stmt_1484/call_stmt_1484_Update/cca
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/EQ_u1_u1_1488_inputs/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/EQ_u1_u1_1488_inputs/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/EQ_u1_u1_1488/SplitProtocol/Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_1415/EQ_u1_u1_1488_place
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_1415/if_stmt_1485_else_link/$entry
      -- 
    cca_1911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1484_call_ack_1, ack => populateRxQueue_CP_1799_elements(12)); -- 
    branch_req_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(12), ack => if_stmt_1485_branch_req_0); -- 
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	21 
    -- CP-element group 13: 	22 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_1415/if_stmt_1485_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_1415/if_stmt_1485_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/$entry
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/$entry
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Sample/req
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Update/req
      -- 
    if_choice_transition_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1485_branch_ack_1, ack => populateRxQueue_CP_1799_elements(13)); -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(13), ack => n_q_index_1475_1427_buf_req_0); -- 
    req_2101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(13), ack => n_q_index_1475_1427_buf_req_1); -- 
    -- CP-element group 14:  merge  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	1 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1415/if_stmt_1485__exit__
      -- CP-element group 14: 	 branch_block_stmt_1415/if_stmt_1485_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_1415/if_stmt_1485_else_link/else_choice_transition
      -- 
    else_choice_transition_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1485_branch_ack_0, ack => populateRxQueue_CP_1799_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Update/req
      -- 
    ack_1962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_ack_0, ack => populateRxQueue_CP_1799_elements(15)); -- 
    req_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(15), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_req_1); -- 
    -- CP-element group 16:  transition  place  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	1 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1415/assign_stmt_1494__exit__
      -- CP-element group 16: 	 branch_block_stmt_1415/assign_stmt_1494/$exit
      -- CP-element group 16: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1415/assign_stmt_1494/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_Update/ack
      -- 
    ack_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_ack_1, ack => populateRxQueue_CP_1799_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (71) 
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Update/req
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/ADD_u6_u6_1421_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/ADD_u6_u6_1421/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Update/req
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SUB_u32_u32_1424_inputs/RPIPE_NUMBER_OF_SERVERS_1422/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SUB_u32_u32_1424/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/AND_u6_u6_1426_inputs/type_cast_1425/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Update/cr
      -- 
    rr_2073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(17), ack => AND_u6_u6_1426_inst_req_0); -- 
    cr_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(17), ack => AND_u6_u6_1426_inst_req_1); -- 
    populateRxQueue_CP_1799_elements(17) <= populateRxQueue_CP_1799_elements(0);
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Sample/ra
      -- 
    ra_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1426_inst_ack_0, ack => populateRxQueue_CP_1799_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/Update/ca
      -- 
    ca_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1426_inst_ack_1, ack => populateRxQueue_CP_1799_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	24 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/$exit
      -- CP-element group 20: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/$exit
      -- CP-element group 20: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/$exit
      -- CP-element group 20: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/$exit
      -- CP-element group 20: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_sources/AND_u6_u6_1426/SplitProtocol/$exit
      -- CP-element group 20: 	 branch_block_stmt_1415/merge_stmt_1416__entry___PhiReq/phi_stmt_1417/phi_stmt_1417_req
      -- 
    phi_stmt_1417_req_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1417_req_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(20), ack => phi_stmt_1417_req_0); -- 
    populateRxQueue_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1799_elements(18) & populateRxQueue_CP_1799_elements(19);
      gj_populateRxQueue_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1799_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	13 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Sample/ack
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1475_1427_buf_ack_0, ack => populateRxQueue_CP_1799_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/Update/ack
      -- 
    ack_2102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1475_1427_buf_ack_1, ack => populateRxQueue_CP_1799_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1415/loopback_PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/$exit
      -- CP-element group 23: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/$exit
      -- CP-element group 23: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_sources/Interlock/$exit
      -- CP-element group 23: 	 branch_block_stmt_1415/loopback_PhiReq/phi_stmt_1417/phi_stmt_1417_req
      -- 
    phi_stmt_1417_req_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1417_req_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(23), ack => phi_stmt_1417_req_1); -- 
    populateRxQueue_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1799_elements(21) & populateRxQueue_CP_1799_elements(22);
      gj_populateRxQueue_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1799_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  merge  transition  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1415/merge_stmt_1416_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_1415/merge_stmt_1416_PhiAck/$entry
      -- 
    populateRxQueue_CP_1799_elements(24) <= OrReduce(populateRxQueue_CP_1799_elements(20) & populateRxQueue_CP_1799_elements(23));
    -- CP-element group 25:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: 	3 
    -- CP-element group 25: 	5 
    -- CP-element group 25: 	6 
    -- CP-element group 25: 	7 
    -- CP-element group 25:  members (20) 
      -- CP-element group 25: 	 branch_block_stmt_1415/merge_stmt_1416__exit__
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475__entry__
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/$entry
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Sample/crr
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1448_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/call_stmt_1465_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1415/assign_stmt_1436_to_assign_stmt_1475/AND_u6_u6_1474_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1415/merge_stmt_1416_PhiAck/$exit
      -- CP-element group 25: 	 branch_block_stmt_1415/merge_stmt_1416_PhiAck/phi_stmt_1417_ack
      -- 
    phi_stmt_1417_ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1417_ack_0, ack => populateRxQueue_CP_1799_elements(25)); -- 
    crr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(25), ack => call_stmt_1448_call_req_0); -- 
    ccr_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(25), ack => call_stmt_1448_call_req_1); -- 
    ccr_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(25), ack => call_stmt_1465_call_req_1); -- 
    rr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(25), ack => AND_u6_u6_1474_inst_req_0); -- 
    cr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1799_elements(25), ack => AND_u6_u6_1474_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1421_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1434_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1469_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_1426_wire : std_logic_vector(5 downto 0);
    signal EQ_u1_u1_1488_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1481_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1443_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1422_wire : std_logic_vector(31 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1470_wire : std_logic_vector(31 downto 0);
    signal R_RX_QUEUES_REG_START_OFFSET_1433_wire_constant : std_logic_vector(5 downto 0);
    signal SUB_u32_u32_1424_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1472_wire : std_logic_vector(31 downto 0);
    signal konst_1420_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1423_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1468_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1471_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1482_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1487_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_1475 : std_logic_vector(5 downto 0);
    signal n_q_index_1475_1427_buffered : std_logic_vector(5 downto 0);
    signal push_status_1465 : std_logic_vector(0 downto 0);
    signal q_index_1417 : std_logic_vector(5 downto 0);
    signal register_index_1436 : std_logic_vector(5 downto 0);
    signal rx_queue_pointer_32_1448 : std_logic_vector(31 downto 0);
    signal rx_queue_pointer_36_1454 : std_logic_vector(35 downto 0);
    signal slice_1463_wire : std_logic_vector(31 downto 0);
    signal status_1484 : std_logic_vector(0 downto 0);
    signal type_cast_1425_wire : std_logic_vector(5 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1451_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1460_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1473_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1443_wire_constant <= "1111";
    R_RX_QUEUES_REG_START_OFFSET_1433_wire_constant <= "000010";
    konst_1420_wire_constant <= "000001";
    konst_1423_wire_constant <= "00000000000000000000000000000001";
    konst_1468_wire_constant <= "000001";
    konst_1471_wire_constant <= "00000000000000000000000000000001";
    konst_1482_wire_constant <= "00000000000000000000000000100000";
    konst_1487_wire_constant <= "0";
    type_cast_1440_wire_constant <= "1";
    type_cast_1446_wire_constant <= "00000000000000000000000000000000";
    type_cast_1451_wire_constant <= "0000";
    type_cast_1460_wire_constant <= "1";
    phi_stmt_1417: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= AND_u6_u6_1426_wire & n_q_index_1475_1427_buffered;
      req <= phi_stmt_1417_req_0 & phi_stmt_1417_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1417",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1417_ack_0,
          idata => idata,
          odata => q_index_1417,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1417
    -- flow-through slice operator slice_1463_inst
    slice_1463_wire <= rx_buffer_pointer_buffer(31 downto 0);
    n_q_index_1475_1427_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_1475_1427_buf_req_0;
      n_q_index_1475_1427_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_1475_1427_buf_req_1;
      n_q_index_1475_1427_buf_ack_1<= rack(0);
      n_q_index_1475_1427_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_1475_1427_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_1475,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_1475_1427_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1425_inst
    process(SUB_u32_u32_1424_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1424_wire(5 downto 0);
      type_cast_1425_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1435_inst
    process(ADD_u6_u6_1434_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1434_wire(5 downto 0);
      register_index_1436 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1473_inst
    process(SUB_u32_u32_1472_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1472_wire(5 downto 0);
      type_cast_1473_wire <= tmp_var; -- 
    end process;
    if_stmt_1479_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1481_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1479_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1479_branch_req_0,
          ack0 => if_stmt_1479_branch_ack_0,
          ack1 => if_stmt_1479_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1485_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_1488_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1485_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1485_branch_req_0,
          ack0 => if_stmt_1485_branch_ack_0,
          ack1 => if_stmt_1485_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u6_u6_1421_inst
    process(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419_wire, konst_1420_wire_constant, tmp_var);
      ADD_u6_u6_1421_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_1434_inst
    process(q_index_1417) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_1417, R_RX_QUEUES_REG_START_OFFSET_1433_wire_constant, tmp_var);
      ADD_u6_u6_1434_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_1469_inst
    process(q_index_1417) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_1417, konst_1468_wire_constant, tmp_var);
      ADD_u6_u6_1469_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_1426_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1421_wire & type_cast_1425_wire;
      AND_u6_u6_1426_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1426_inst_req_0;
      AND_u6_u6_1426_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1426_inst_req_1;
      AND_u6_u6_1426_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : AND_u6_u6_1474_inst 
    ApIntAnd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1469_wire & type_cast_1473_wire;
      n_q_index_1475 <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1474_inst_req_0;
      AND_u6_u6_1474_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1474_inst_req_1;
      AND_u6_u6_1474_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator CONCAT_u4_u36_1453_inst
    process(type_cast_1451_wire_constant, rx_queue_pointer_32_1448) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1451_wire_constant, rx_queue_pointer_32_1448, tmp_var);
      rx_queue_pointer_36_1454 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1488_inst
    process(status_1484) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_1484, konst_1487_wire_constant, tmp_var);
      EQ_u1_u1_1488_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1481_inst
    process(push_status_1465) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_1465, tmp_var);
      NOT_u1_u1_1481_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u32_u32_1424_inst
    process(RPIPE_NUMBER_OF_SERVERS_1422_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1422_wire, konst_1423_wire_constant, tmp_var);
      SUB_u32_u32_1424_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1472_inst
    process(RPIPE_NUMBER_OF_SERVERS_1470_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1470_wire, konst_1471_wire_constant, tmp_var);
      SUB_u32_u32_1472_wire <= tmp_var; --
    end process;
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1419_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_1470_wire <= NUMBER_OF_SERVERS;
    RPIPE_NUMBER_OF_SERVERS_1422_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1492_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_1417;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1448_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1448_call_req_0;
      call_stmt_1448_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1448_call_req_1;
      call_stmt_1448_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1440_wire_constant & NOT_u4_u4_1443_wire_constant & register_index_1436 & type_cast_1446_wire_constant;
      rx_queue_pointer_32_1448 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1465_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1465_call_req_0;
      call_stmt_1465_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1465_call_req_1;
      call_stmt_1465_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1460_wire_constant & rx_queue_pointer_36_1454 & slice_1463_wire;
      push_status_1465 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    operator_delay_time_3273_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_1484_call_req_0;
      call_stmt_1484_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_1484_call_req_1;
      call_stmt_1484_call_ack_1<= update_ack(0);
      call_stmt_1484_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_1482_wire_constant,
        delay_done => status_1484,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(35 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(35 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
    updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(35 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(99 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 69)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_1548_start: Boolean;
  signal pushIntoQueue_CP_1548_symbol: Boolean;
  -- volatile/operator module components. 
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1319_call_ack_0 : boolean;
  signal NOT_u1_u1_1383_inst_req_1 : boolean;
  signal call_stmt_1376_call_ack_0 : boolean;
  signal call_stmt_1319_call_ack_1 : boolean;
  signal call_stmt_1376_call_req_0 : boolean;
  signal call_stmt_1330_call_req_1 : boolean;
  signal call_stmt_1330_call_ack_1 : boolean;
  signal call_stmt_1319_call_req_0 : boolean;
  signal call_stmt_1305_call_req_1 : boolean;
  signal call_stmt_1369_call_ack_1 : boolean;
  signal call_stmt_1305_call_ack_1 : boolean;
  signal call_stmt_1330_call_ack_0 : boolean;
  signal call_stmt_1330_call_req_0 : boolean;
  signal call_stmt_1376_call_req_1 : boolean;
  signal call_stmt_1376_call_ack_1 : boolean;
  signal call_stmt_1364_call_ack_0 : boolean;
  signal NOT_u1_u1_1383_inst_req_0 : boolean;
  signal call_stmt_1319_call_req_1 : boolean;
  signal call_stmt_1364_call_req_0 : boolean;
  signal call_stmt_1333_call_req_0 : boolean;
  signal call_stmt_1333_call_ack_0 : boolean;
  signal NOT_u1_u1_1383_inst_ack_0 : boolean;
  signal call_stmt_1369_call_req_1 : boolean;
  signal call_stmt_1380_call_ack_1 : boolean;
  signal call_stmt_1380_call_req_1 : boolean;
  signal call_stmt_1327_call_ack_1 : boolean;
  signal call_stmt_1327_call_req_1 : boolean;
  signal call_stmt_1369_call_ack_0 : boolean;
  signal call_stmt_1369_call_req_0 : boolean;
  signal NOT_u1_u1_1383_inst_ack_1 : boolean;
  signal call_stmt_1305_call_ack_0 : boolean;
  signal call_stmt_1333_call_ack_1 : boolean;
  signal call_stmt_1305_call_req_0 : boolean;
  signal call_stmt_1380_call_ack_0 : boolean;
  signal call_stmt_1380_call_req_0 : boolean;
  signal call_stmt_1327_call_ack_0 : boolean;
  signal call_stmt_1327_call_req_0 : boolean;
  signal call_stmt_1333_call_req_1 : boolean;
  signal call_stmt_1364_call_ack_1 : boolean;
  signal call_stmt_1364_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 69) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(68 downto 37) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(68 downto 37);
  in_buffer_data_in(tag_length + 68 downto 69) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 68 downto 69);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_1548_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1548_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1548_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1548_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_1548: Block -- control-path 
    signal pushIntoQueue_CP_1548_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_1548_elements(0) <= pushIntoQueue_CP_1548_start;
    pushIntoQueue_CP_1548_symbol <= pushIntoQueue_CP_1548_elements(24);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_update_start_
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Update/$entry
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_update_start_
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_sample_start_
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Update/ccr
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Update/ccr
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Update/$entry
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Sample/crr
      -- CP-element group 0: 	 call_stmt_1305_to_call_stmt_1319/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(0), ack => call_stmt_1305_call_req_0); -- 
    ccr_1566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(0), ack => call_stmt_1305_call_req_1); -- 
    ccr_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(0), ack => call_stmt_1319_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_sample_completed_
      -- CP-element group 1: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Sample/cra
      -- 
    cra_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1305_call_ack_0, ack => pushIntoQueue_CP_1548_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Sample/crr
      -- CP-element group 2: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Update/cca
      -- CP-element group 2: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_update_completed_
      -- CP-element group 2: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_sample_start_
      -- CP-element group 2: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1305_Update/$exit
      -- 
    cca_1567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1305_call_ack_1, ack => pushIntoQueue_CP_1548_elements(2)); -- 
    crr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(2), ack => call_stmt_1319_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Sample/cra
      -- CP-element group 3: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_sample_completed_
      -- CP-element group 3: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Sample/$exit
      -- 
    cra_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1319_call_ack_0, ack => pushIntoQueue_CP_1548_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	16 
    -- CP-element group 4: 	19 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	13 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	8 
    -- CP-element group 4:  members (26) 
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/$entry
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Update/$entry
      -- CP-element group 4: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Update/cca
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_update_start_
      -- CP-element group 4: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_update_completed_
      -- CP-element group 4: 	 call_stmt_1305_to_call_stmt_1319/$exit
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Update/ccr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Update/$entry
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Update/ccr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_sample_start_
      -- CP-element group 4: 	 call_stmt_1305_to_call_stmt_1319/call_stmt_1319_Update/$exit
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_update_start_
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_update_start_
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_update_start_
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Update/$entry
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Update/ccr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Update/$entry
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_update_start_
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Update/ccr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Update/$entry
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Sample/crr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_update_start_
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Update/ccr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Update/ccr
      -- CP-element group 4: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Update/$entry
      -- 
    cca_1581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1319_call_ack_1, ack => pushIntoQueue_CP_1548_elements(4)); -- 
    ccr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1376_call_req_1); -- 
    ccr_1625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1333_call_req_1); -- 
    ccr_1639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1364_call_req_1); -- 
    ccr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1369_call_req_1); -- 
    crr_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1327_call_req_0); -- 
    ccr_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1327_call_req_1); -- 
    ccr_1611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(4), ack => call_stmt_1330_call_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_sample_completed_
      -- CP-element group 5: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Sample/cra
      -- CP-element group 5: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Sample/$exit
      -- 
    cra_1593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1327_call_ack_0, ack => pushIntoQueue_CP_1548_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	17 
    -- CP-element group 6: 	11 
    -- CP-element group 6: 	14 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Sample/crr
      -- CP-element group 6: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_update_completed_
      -- CP-element group 6: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_sample_start_
      -- CP-element group 6: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Update/cca
      -- CP-element group 6: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1327_Update/$exit
      -- 
    cca_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1327_call_ack_1, ack => pushIntoQueue_CP_1548_elements(6)); -- 
    crr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(6), ack => call_stmt_1330_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Sample/cra
      -- CP-element group 7: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Sample/$exit
      -- CP-element group 7: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_sample_completed_
      -- 
    cra_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1330_call_ack_0, ack => pushIntoQueue_CP_1548_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	17 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_sample_start_
      -- CP-element group 8: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Update/cca
      -- CP-element group 8: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_Update/$exit
      -- CP-element group 8: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Sample/crr
      -- CP-element group 8: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1330_update_completed_
      -- 
    cca_1612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1330_call_ack_1, ack => pushIntoQueue_CP_1548_elements(8)); -- 
    crr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(8), ack => call_stmt_1333_call_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Sample/$exit
      -- CP-element group 9: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_sample_completed_
      -- CP-element group 9: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Sample/cra
      -- 
    cra_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1333_call_ack_0, ack => pushIntoQueue_CP_1548_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_update_completed_
      -- CP-element group 10: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Update/$exit
      -- CP-element group 10: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1333_Update/cca
      -- 
    cca_1626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1333_call_ack_1, ack => pushIntoQueue_CP_1548_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_sample_start_
      -- CP-element group 11: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Sample/$entry
      -- CP-element group 11: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Sample/crr
      -- 
    crr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(11), ack => call_stmt_1364_call_req_0); -- 
    pushIntoQueue_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1548_elements(10) & pushIntoQueue_CP_1548_elements(6) & pushIntoQueue_CP_1548_elements(8);
      gj_pushIntoQueue_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1548_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_sample_completed_
      -- CP-element group 12: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Sample/$exit
      -- CP-element group 12: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Sample/cra
      -- 
    cra_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1364_call_ack_0, ack => pushIntoQueue_CP_1548_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	4 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_update_completed_
      -- CP-element group 13: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Update/cca
      -- CP-element group 13: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1364_Update/$exit
      -- 
    cca_1640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1364_call_ack_1, ack => pushIntoQueue_CP_1548_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: 	6 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Sample/crr
      -- CP-element group 14: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Sample/$entry
      -- CP-element group 14: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_sample_start_
      -- 
    crr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(14), ack => call_stmt_1369_call_req_0); -- 
    pushIntoQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1548_elements(13) & pushIntoQueue_CP_1548_elements(6) & pushIntoQueue_CP_1548_elements(8);
      gj_pushIntoQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1548_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Sample/cra
      -- CP-element group 15: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Sample/$exit
      -- CP-element group 15: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_sample_completed_
      -- 
    cra_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1369_call_ack_0, ack => pushIntoQueue_CP_1548_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	4 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Update/cca
      -- CP-element group 16: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_Update/$exit
      -- CP-element group 16: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1369_update_completed_
      -- 
    cca_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1369_call_ack_1, ack => pushIntoQueue_CP_1548_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: 	10 
    -- CP-element group 17: 	6 
    -- CP-element group 17: 	8 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Sample/$entry
      -- CP-element group 17: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Sample/crr
      -- CP-element group 17: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_sample_start_
      -- 
    crr_1662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(17), ack => call_stmt_1376_call_req_0); -- 
    pushIntoQueue_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1548_elements(16) & pushIntoQueue_CP_1548_elements(10) & pushIntoQueue_CP_1548_elements(6) & pushIntoQueue_CP_1548_elements(8);
      gj_pushIntoQueue_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1548_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Sample/cra
      -- CP-element group 18: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_sample_completed_
      -- 
    cra_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1376_call_ack_0, ack => pushIntoQueue_CP_1548_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (17) 
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Update/cr
      -- CP-element group 19: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_update_completed_
      -- CP-element group 19: 	 call_stmt_1327_to_call_stmt_1376/$exit
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/$entry
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_update_start_
      -- CP-element group 19: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Update/$exit
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_sample_start_
      -- CP-element group 19: 	 call_stmt_1327_to_call_stmt_1376/call_stmt_1376_Update/cca
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Sample/rr
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Update/$entry
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Update/ccr
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Update/$entry
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Sample/crr
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_update_start_
      -- CP-element group 19: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_sample_start_
      -- 
    cca_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1376_call_ack_1, ack => pushIntoQueue_CP_1548_elements(19)); -- 
    crr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(19), ack => call_stmt_1380_call_req_0); -- 
    ccr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(19), ack => call_stmt_1380_call_req_1); -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(19), ack => NOT_u1_u1_1383_inst_req_0); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1548_elements(19), ack => NOT_u1_u1_1383_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Sample/cra
      -- CP-element group 20: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_sample_completed_
      -- 
    cra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1380_call_ack_0, ack => pushIntoQueue_CP_1548_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Update/cca
      -- CP-element group 21: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_Update/$exit
      -- CP-element group 21: 	 call_stmt_1380_to_assign_stmt_1384/call_stmt_1380_update_completed_
      -- 
    cca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1380_call_ack_1, ack => pushIntoQueue_CP_1548_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Sample/$exit
      -- CP-element group 22: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_sample_completed_
      -- CP-element group 22: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Sample/ra
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1383_inst_ack_0, ack => pushIntoQueue_CP_1548_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Update/$exit
      -- CP-element group 23: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_update_completed_
      -- CP-element group 23: 	 call_stmt_1380_to_assign_stmt_1384/NOT_u1_u1_1383_Update/ca
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1383_inst_ack_1, ack => pushIntoQueue_CP_1548_elements(23)); -- 
    -- CP-element group 24:  join  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 $exit
      -- CP-element group 24: 	 call_stmt_1380_to_assign_stmt_1384/$exit
      -- 
    pushIntoQueue_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1548_elements(21) & pushIntoQueue_CP_1548_elements(23);
      gj_pushIntoQueue_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1548_elements(24), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1346_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1375_wire : std_logic_vector(31 downto 0);
    signal ADD_u36_u36_1301_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_1298_wire_constant : std_logic_vector(7 downto 0);
    signal Queue_Length_1330 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1338_wire : std_logic_vector(31 downto 0);
    signal ba_and_misc_1305 : std_logic_vector(63 downto 0);
    signal konst_1300_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1337_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1343_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1345_wire_constant : std_logic_vector(31 downto 0);
    signal lock_n_1315 : std_logic_vector(0 downto 0);
    signal m_ok_1319 : std_logic_vector(0 downto 0);
    signal misc_1309 : std_logic_vector(31 downto 0);
    signal next_wi_1348 : std_logic_vector(31 downto 0);
    signal q_full_1353 : std_logic_vector(0 downto 0);
    signal read_index_1327 : std_logic_vector(31 downto 0);
    signal round_off_1340 : std_logic_vector(0 downto 0);
    signal total_msgs_1333 : std_logic_vector(31 downto 0);
    signal type_cast_1293_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1295_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1303_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1313_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1374_wire_constant : std_logic_vector(31 downto 0);
    signal write_index_1327 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_1298_wire_constant <= "11111111";
    konst_1300_wire_constant <= "000000000000000000000000000000011000";
    konst_1337_wire_constant <= "00000000000000000000000000000001";
    konst_1343_wire_constant <= "00000000000000000000000000000000";
    konst_1345_wire_constant <= "00000000000000000000000000000001";
    type_cast_1293_wire_constant <= "0";
    type_cast_1295_wire_constant <= "1";
    type_cast_1303_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1313_wire_constant <= "00000000000000000000000000000000";
    type_cast_1374_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_1347_inst
    next_wi_1348 <= konst_1343_wire_constant when (round_off_1340(0) /=  '0') else ADD_u32_u32_1346_wire;
    -- flow-through slice operator slice_1308_inst
    misc_1309 <= ba_and_misc_1305(31 downto 0);
    -- binary operator ADD_u32_u32_1346_inst
    process(write_index_1327) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(write_index_1327, konst_1345_wire_constant, tmp_var);
      ADD_u32_u32_1346_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1375_inst
    process(total_msgs_1333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(total_msgs_1333, type_cast_1374_wire_constant, tmp_var);
      ADD_u32_u32_1375_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_1301_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_1300_wire_constant, tmp_var);
      ADD_u36_u36_1301_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1314_inst
    process(misc_1309) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(misc_1309, type_cast_1313_wire_constant, tmp_var);
      lock_n_1315 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1339_inst
    process(write_index_1327, SUB_u32_u32_1338_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_1327, SUB_u32_u32_1338_wire, tmp_var);
      round_off_1340 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1352_inst
    process(next_wi_1348, read_index_1327) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_wi_1348, read_index_1327, tmp_var);
      q_full_1353 <= tmp_var; --
    end process;
    -- shared split operator group (6) : NOT_u1_u1_1383_inst 
    ApIntNot_group_6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_full_1353;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1383_inst_req_0;
      NOT_u1_u1_1383_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1383_inst_req_1;
      NOT_u1_u1_1383_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_6_gI: SplitGuardInterface generic map(name => "ApIntNot_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- binary operator SUB_u32_u32_1338_inst
    process(Queue_Length_1330) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(Queue_Length_1330, konst_1337_wire_constant, tmp_var);
      SUB_u32_u32_1338_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1305_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1305_call_req_0;
      call_stmt_1305_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1305_call_req_1;
      call_stmt_1305_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1293_wire_constant & type_cast_1295_wire_constant & NOT_u8_u8_1298_wire_constant & ADD_u36_u36_1301_wire & type_cast_1303_wire_constant;
      ba_and_misc_1305 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1319_call 
    acquireLock_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1319_call_req_0;
      call_stmt_1319_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1319_call_req_1;
      call_stmt_1319_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_1315(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_1_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_1319 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(35 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1327_call 
    getQueuePointers_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1327_call_req_0;
      call_stmt_1327_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1327_call_req_1;
      call_stmt_1327_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_2_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_index_1327 <= data_out(63 downto 32);
      read_index_1327 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1330_call 
    getQueueLength_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1330_call_req_0;
      call_stmt_1330_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1330_call_req_1;
      call_stmt_1330_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_3_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      Queue_Length_1330 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(35 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1333_call 
    getTotalMessages_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1333_call_req_0;
      call_stmt_1333_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1333_call_req_1;
      call_stmt_1333_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_4_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      total_msgs_1333 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(35 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1364_call 
    setQueueElement_call_group_5: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1364_call_req_0;
      call_stmt_1364_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1364_call_req_1;
      call_stmt_1364_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1353(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_5_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_index_1327 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(99 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1369_call 
    setQueuePointers_call_group_6: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1369_call_req_0;
      call_stmt_1369_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1369_call_req_1;
      call_stmt_1369_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1353(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_6_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & next_wi_1348 & read_index_1327;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1376_call 
    updateTotalMessages_call_group_7: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1376_call_req_0;
      call_stmt_1376_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1376_call_req_1;
      call_stmt_1376_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1353(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateTotalMessages_call_group_7_gI: SplitGuardInterface generic map(name => "updateTotalMessages_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & ADD_u32_u32_1375_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateTotalMessages_call_reqs(0),
          ackR => updateTotalMessages_call_acks(0),
          dataR => updateTotalMessages_call_data(67 downto 0),
          tagR => updateTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => updateTotalMessages_return_acks(0), -- cross-over
          ackL => updateTotalMessages_return_reqs(0), -- cross-over
          tagL => updateTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_1380_call 
    releaseLock_call_group_8: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1380_call_req_0;
      call_stmt_1380_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1380_call_req_1;
      call_stmt_1380_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_1315(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_8_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(35 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity releaseLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseLock;
architecture releaseLock_arch of releaseLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal releaseLock_CP_910_start: Boolean;
  signal releaseLock_CP_910_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_935_call_ack_0 : boolean;
  signal call_stmt_935_call_ack_1 : boolean;
  signal call_stmt_935_call_req_1 : boolean;
  signal call_stmt_817_call_req_1 : boolean;
  signal call_stmt_817_call_req_0 : boolean;
  signal call_stmt_935_call_req_0 : boolean;
  signal call_stmt_817_call_ack_0 : boolean;
  signal call_stmt_817_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseLock_CP_910_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_910_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseLock_CP_910_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_910_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseLock_CP_910: Block -- control-path 
    signal releaseLock_CP_910_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    releaseLock_CP_910_elements(0) <= releaseLock_CP_910_start;
    releaseLock_CP_910_symbol <= releaseLock_CP_910_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_update_start_
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Update/ccr
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Update/ccr
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Sample/crr
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Update/$entry
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Update/$entry
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_sample_start_
      -- CP-element group 0: 	 assign_stmt_805_to_call_stmt_935/$entry
      -- 
    crr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_910_elements(0), ack => call_stmt_817_call_req_0); -- 
    ccr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_910_elements(0), ack => call_stmt_817_call_req_1); -- 
    ccr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_910_elements(0), ack => call_stmt_935_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_sample_completed_
      -- CP-element group 1: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Sample/cra
      -- 
    cra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_817_call_ack_0, ack => releaseLock_CP_910_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_update_completed_
      -- CP-element group 2: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_sample_start_
      -- CP-element group 2: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Sample/crr
      -- CP-element group 2: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Update/$exit
      -- CP-element group 2: 	 assign_stmt_805_to_call_stmt_935/call_stmt_817_Update/cca
      -- 
    cca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_817_call_ack_1, ack => releaseLock_CP_910_elements(2)); -- 
    crr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_910_elements(2), ack => call_stmt_935_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Sample/cra
      -- CP-element group 3: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_sample_completed_
      -- CP-element group 3: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Sample/$exit
      -- 
    cra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_935_call_ack_0, ack => releaseLock_CP_910_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Update/cca
      -- CP-element group 4: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_Update/$exit
      -- CP-element group 4: 	 assign_stmt_805_to_call_stmt_935/call_stmt_935_update_completed_
      -- CP-element group 4: 	 assign_stmt_805_to_call_stmt_935/$exit
      -- CP-element group 4: 	 $exit
      -- 
    cca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_935_call_ack_1, ack => releaseLock_CP_910_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_879_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_892_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_906_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_919_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_893_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_920_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u4_u36_931_wire : std_logic_vector(35 downto 0);
    signal MUX_872_wire : std_logic_vector(0 downto 0);
    signal MUX_878_wire : std_logic_vector(0 downto 0);
    signal MUX_885_wire : std_logic_vector(0 downto 0);
    signal MUX_891_wire : std_logic_vector(0 downto 0);
    signal MUX_899_wire : std_logic_vector(0 downto 0);
    signal MUX_905_wire : std_logic_vector(0 downto 0);
    signal MUX_912_wire : std_logic_vector(0 downto 0);
    signal MUX_918_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_812_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_935 : std_logic_vector(63 downto 0);
    signal konst_828_wire_constant : std_logic_vector(2 downto 0);
    signal konst_833_wire_constant : std_logic_vector(2 downto 0);
    signal konst_838_wire_constant : std_logic_vector(2 downto 0);
    signal konst_843_wire_constant : std_logic_vector(2 downto 0);
    signal konst_848_wire_constant : std_logic_vector(2 downto 0);
    signal konst_853_wire_constant : std_logic_vector(2 downto 0);
    signal konst_858_wire_constant : std_logic_vector(2 downto 0);
    signal konst_863_wire_constant : std_logic_vector(2 downto 0);
    signal lock_addr_32_821 : std_logic_vector(31 downto 0);
    signal lock_address_pointer_805 : std_logic_vector(35 downto 0);
    signal msg_size_plus_lock_817 : std_logic_vector(63 downto 0);
    signal new_bmask_922 : std_logic_vector(7 downto 0);
    signal s0_830 : std_logic_vector(0 downto 0);
    signal s1_835 : std_logic_vector(0 downto 0);
    signal s2_840 : std_logic_vector(0 downto 0);
    signal s3_845 : std_logic_vector(0 downto 0);
    signal s4_850 : std_logic_vector(0 downto 0);
    signal s5_855 : std_logic_vector(0 downto 0);
    signal s6_860 : std_logic_vector(0 downto 0);
    signal s7_865 : std_logic_vector(0 downto 0);
    signal sel_825 : std_logic_vector(2 downto 0);
    signal type_cast_803_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_807_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_815_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_869_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_871_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_875_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_877_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_882_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_884_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_888_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_896_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_902_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_904_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_909_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_911_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_917_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_924_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_929_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_933_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_812_wire_constant <= "11111111";
    konst_828_wire_constant <= "000";
    konst_833_wire_constant <= "001";
    konst_838_wire_constant <= "010";
    konst_843_wire_constant <= "011";
    konst_848_wire_constant <= "100";
    konst_853_wire_constant <= "101";
    konst_858_wire_constant <= "110";
    konst_863_wire_constant <= "111";
    type_cast_803_wire_constant <= "000000000000000000000000000000010000";
    type_cast_807_wire_constant <= "1";
    type_cast_809_wire_constant <= "1";
    type_cast_815_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_869_wire_constant <= "1";
    type_cast_871_wire_constant <= "0";
    type_cast_875_wire_constant <= "1";
    type_cast_877_wire_constant <= "0";
    type_cast_882_wire_constant <= "1";
    type_cast_884_wire_constant <= "0";
    type_cast_888_wire_constant <= "1";
    type_cast_890_wire_constant <= "0";
    type_cast_896_wire_constant <= "1";
    type_cast_898_wire_constant <= "0";
    type_cast_902_wire_constant <= "1";
    type_cast_904_wire_constant <= "0";
    type_cast_909_wire_constant <= "1";
    type_cast_911_wire_constant <= "0";
    type_cast_915_wire_constant <= "1";
    type_cast_917_wire_constant <= "0";
    type_cast_924_wire_constant <= "0";
    type_cast_926_wire_constant <= "0";
    type_cast_929_wire_constant <= "0000";
    type_cast_933_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_872_inst
    MUX_872_wire <= type_cast_869_wire_constant when (s0_830(0) /=  '0') else type_cast_871_wire_constant;
    -- flow-through select operator MUX_878_inst
    MUX_878_wire <= type_cast_875_wire_constant when (s1_835(0) /=  '0') else type_cast_877_wire_constant;
    -- flow-through select operator MUX_885_inst
    MUX_885_wire <= type_cast_882_wire_constant when (s2_840(0) /=  '0') else type_cast_884_wire_constant;
    -- flow-through select operator MUX_891_inst
    MUX_891_wire <= type_cast_888_wire_constant when (s3_845(0) /=  '0') else type_cast_890_wire_constant;
    -- flow-through select operator MUX_899_inst
    MUX_899_wire <= type_cast_896_wire_constant when (s4_850(0) /=  '0') else type_cast_898_wire_constant;
    -- flow-through select operator MUX_905_inst
    MUX_905_wire <= type_cast_902_wire_constant when (s5_855(0) /=  '0') else type_cast_904_wire_constant;
    -- flow-through select operator MUX_912_inst
    MUX_912_wire <= type_cast_909_wire_constant when (s6_860(0) /=  '0') else type_cast_911_wire_constant;
    -- flow-through select operator MUX_918_inst
    MUX_918_wire <= type_cast_915_wire_constant when (s7_865(0) /=  '0') else type_cast_917_wire_constant;
    -- flow-through slice operator slice_820_inst
    lock_addr_32_821 <= msg_size_plus_lock_817(31 downto 0);
    -- flow-through slice operator slice_824_inst
    sel_825 <= lock_addr_32_821(2 downto 0);
    -- binary operator ADD_u36_u36_804_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_803_wire_constant, tmp_var);
      lock_address_pointer_805 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_879_inst
    process(MUX_872_wire, MUX_878_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_872_wire, MUX_878_wire, tmp_var);
      CONCAT_u1_u2_879_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_892_inst
    process(MUX_885_wire, MUX_891_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_885_wire, MUX_891_wire, tmp_var);
      CONCAT_u1_u2_892_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_906_inst
    process(MUX_899_wire, MUX_905_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_899_wire, MUX_905_wire, tmp_var);
      CONCAT_u1_u2_906_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_919_inst
    process(MUX_912_wire, MUX_918_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_912_wire, MUX_918_wire, tmp_var);
      CONCAT_u1_u2_919_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_893_inst
    process(CONCAT_u1_u2_879_wire, CONCAT_u1_u2_892_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_879_wire, CONCAT_u1_u2_892_wire, tmp_var);
      CONCAT_u2_u4_893_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_920_inst
    process(CONCAT_u1_u2_906_wire, CONCAT_u1_u2_919_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_906_wire, CONCAT_u1_u2_919_wire, tmp_var);
      CONCAT_u2_u4_920_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_931_inst
    process(type_cast_929_wire_constant, lock_addr_32_821) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_929_wire_constant, lock_addr_32_821, tmp_var);
      CONCAT_u4_u36_931_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_921_inst
    process(CONCAT_u2_u4_893_wire, CONCAT_u2_u4_920_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_893_wire, CONCAT_u2_u4_920_wire, tmp_var);
      new_bmask_922 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_829_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_828_wire_constant, tmp_var);
      s0_830 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_834_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_833_wire_constant, tmp_var);
      s1_835 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_839_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_838_wire_constant, tmp_var);
      s2_840 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_844_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_843_wire_constant, tmp_var);
      s3_845 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_849_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_848_wire_constant, tmp_var);
      s4_850 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_854_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_853_wire_constant, tmp_var);
      s5_855 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_859_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_858_wire_constant, tmp_var);
      s6_860 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_864_inst
    process(sel_825) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_825, konst_863_wire_constant, tmp_var);
      s7_865 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_817_call call_stmt_935_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_817_call_req_0;
      reqL_unguarded(0) <= call_stmt_935_call_req_0;
      call_stmt_817_call_ack_0 <= ackL_unguarded(1);
      call_stmt_935_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_817_call_req_1;
      reqR_unguarded(0) <= call_stmt_935_call_req_1;
      call_stmt_817_call_ack_1 <= ackR_unguarded(1);
      call_stmt_935_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_807_wire_constant & type_cast_809_wire_constant & NOT_u8_u8_812_wire_constant & lock_address_pointer_805 & type_cast_815_wire_constant & type_cast_924_wire_constant & type_cast_926_wire_constant & new_bmask_922 & CONCAT_u4_u36_931_wire & type_cast_933_wire_constant;
      msg_size_plus_lock_817 <= data_out(127 downto 64);
      ignore_935 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    write_index : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal write_index_buffer :  std_logic_vector(31 downto 0);
  signal write_index_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_1528_start: Boolean;
  signal setQueueElement_CP_1528_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1285_call_req_0 : boolean;
  signal call_stmt_1285_call_ack_1 : boolean;
  signal call_stmt_1285_call_req_1 : boolean;
  signal call_stmt_1285_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= write_index;
  write_index_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_1528_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1528_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_1528_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1528_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_1528: Block -- control-path 
    signal setQueueElement_CP_1528_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_1528_elements(0) <= setQueueElement_CP_1528_start;
    setQueueElement_CP_1528_symbol <= setQueueElement_CP_1528_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_update_start_
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/$entry
      -- CP-element group 0: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_sample_start_
      -- CP-element group 0: 	 $entry
      -- 
    ccr_1546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1528_elements(0), ack => call_stmt_1285_call_req_1); -- 
    crr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1528_elements(0), ack => call_stmt_1285_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Sample/cra
      -- 
    cra_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1285_call_ack_0, ack => setQueueElement_CP_1528_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_update_completed_
      -- CP-element group 2: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Update/cca
      -- CP-element group 2: 	 assign_stmt_1229_to_call_stmt_1285/$exit
      -- CP-element group 2: 	 assign_stmt_1229_to_call_stmt_1285/call_stmt_1285_Update/$exit
      -- CP-element group 2: 	 $exit
      -- 
    cca_1547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1285_call_ack_1, ack => setQueueElement_CP_1528_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1243_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1261_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_1236_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u32_u64_1265_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1269_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_1249_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_1255_wire_constant : std_logic_vector(7 downto 0);
    signal bmask_1257 : std_logic_vector(7 downto 0);
    signal buffer_address_1229 : std_logic_vector(35 downto 0);
    signal element_pair_address_1239 : std_logic_vector(35 downto 0);
    signal ignore_1285 : std_logic_vector(63 downto 0);
    signal konst_1242_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1260_wire_constant : std_logic_vector(31 downto 0);
    signal slice_1233_wire : std_logic_vector(30 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_1235_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1237_wire : std_logic_vector(35 downto 0);
    signal type_cast_1263_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1278_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1280_wire_constant : std_logic_vector(0 downto 0);
    signal wval_1271 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_1249_wire_constant <= "00001111";
    CONCAT_u4_u8_1255_wire_constant <= "11110000";
    konst_1242_wire_constant <= "00000000000000000000000000000000";
    konst_1260_wire_constant <= "00000000000000000000000000000000";
    type_cast_1227_wire_constant <= "000000000000000000000000000000100000";
    type_cast_1235_wire_constant <= "000";
    type_cast_1263_wire_constant <= "00000000000000000000000000000000";
    type_cast_1268_wire_constant <= "00000000000000000000000000000000";
    type_cast_1278_wire_constant <= "0";
    type_cast_1280_wire_constant <= "0";
    -- flow-through select operator MUX_1256_inst
    bmask_1257 <= CONCAT_u4_u8_1249_wire_constant when (BITSEL_u32_u1_1243_wire(0) /=  '0') else CONCAT_u4_u8_1255_wire_constant;
    -- flow-through select operator MUX_1270_inst
    wval_1271 <= CONCAT_u32_u64_1265_wire when (BITSEL_u32_u1_1261_wire(0) /=  '0') else CONCAT_u32_u64_1269_wire;
    -- flow-through slice operator slice_1233_inst
    slice_1233_wire <= write_index_buffer(31 downto 1);
    -- interlock type_cast_1237_inst
    process(CONCAT_u31_u34_1236_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_1236_wire(33 downto 0);
      type_cast_1237_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_1228_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_1227_wire_constant, tmp_var);
      buffer_address_1229 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_1238_inst
    process(buffer_address_1229, type_cast_1237_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_1229, type_cast_1237_wire, tmp_var);
      element_pair_address_1239 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1243_inst
    process(write_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_index_buffer, konst_1242_wire_constant, tmp_var);
      BITSEL_u32_u1_1243_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1261_inst
    process(write_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_index_buffer, konst_1260_wire_constant, tmp_var);
      BITSEL_u32_u1_1261_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_1236_inst
    process(slice_1233_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1233_wire, type_cast_1235_wire_constant, tmp_var);
      CONCAT_u31_u34_1236_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_1265_inst
    process(type_cast_1263_wire_constant, q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1263_wire_constant, q_w_data_buffer, tmp_var);
      CONCAT_u32_u64_1265_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_1269_inst
    process(q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(q_w_data_buffer, type_cast_1268_wire_constant, tmp_var);
      CONCAT_u32_u64_1269_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1285_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1285_call_req_0;
      call_stmt_1285_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1285_call_req_1;
      call_stmt_1285_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1278_wire_constant & type_cast_1280_wire_constant & bmask_1257 & element_pair_address_1239 & wval_1271;
      ignore_1285 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_856_start: Boolean;
  signal setQueuePointers_CP_856_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_776_call_req_1 : boolean;
  signal call_stmt_758_call_req_1 : boolean;
  signal call_stmt_758_call_ack_1 : boolean;
  signal call_stmt_758_call_req_0 : boolean;
  signal call_stmt_776_call_ack_1 : boolean;
  signal call_stmt_758_call_ack_0 : boolean;
  signal call_stmt_776_call_ack_0 : boolean;
  signal call_stmt_776_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= wp;
  wp_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= rp;
  rp_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_856_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_856_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_856_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_856_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_856: Block -- control-path 
    signal setQueuePointers_CP_856_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_856_elements(0) <= setQueuePointers_CP_856_start;
    setQueuePointers_CP_856_symbol <= setQueuePointers_CP_856_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_sample_start_
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Update/$entry
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Sample/$entry
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Update/ccr
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Update/ccr
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_update_start_
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Sample/crr
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Update/$entry
      -- CP-element group 0: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_update_start_
      -- 
    crr_869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_856_elements(0), ack => call_stmt_758_call_req_0); -- 
    ccr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_856_elements(0), ack => call_stmt_758_call_req_1); -- 
    ccr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_856_elements(0), ack => call_stmt_776_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_sample_completed_
      -- CP-element group 1: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Sample/$exit
      -- CP-element group 1: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Sample/cra
      -- 
    cra_870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_758_call_ack_0, ack => setQueuePointers_CP_856_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_update_completed_
      -- CP-element group 2: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Update/$exit
      -- CP-element group 2: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_sample_start_
      -- CP-element group 2: 	 call_stmt_758_to_call_stmt_776/call_stmt_758_Update/cca
      -- CP-element group 2: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Sample/crr
      -- CP-element group 2: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Sample/$entry
      -- 
    cca_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_758_call_ack_1, ack => setQueuePointers_CP_856_elements(2)); -- 
    crr_883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_856_elements(2), ack => call_stmt_776_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_sample_completed_
      -- CP-element group 3: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Sample/cra
      -- CP-element group 3: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Sample/$exit
      -- 
    cra_884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_776_call_ack_0, ack => setQueuePointers_CP_856_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Update/$exit
      -- CP-element group 4: 	 call_stmt_758_to_call_stmt_776/$exit
      -- CP-element group 4: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_Update/cca
      -- CP-element group 4: 	 call_stmt_758_to_call_stmt_776/call_stmt_776_update_completed_
      -- 
    cca_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_776_call_ack_1, ack => setQueuePointers_CP_856_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_771_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u32_u64_756_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_774_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_752_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_768_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_1_776 : std_logic_vector(63 downto 0);
    signal ignore_758 : std_logic_vector(63 downto 0);
    signal konst_770_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_744_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_762_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_752_wire_constant <= "00001111";
    CONCAT_u4_u8_768_wire_constant <= "11110000";
    konst_770_wire_constant <= "000000000000000000000000000000001000";
    type_cast_744_wire_constant <= "0";
    type_cast_746_wire_constant <= "0";
    type_cast_760_wire_constant <= "0";
    type_cast_762_wire_constant <= "0";
    -- binary operator ADD_u36_u36_771_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_770_wire_constant, tmp_var);
      ADD_u36_u36_771_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_756_inst
    process(rp_buffer, rp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(rp_buffer, rp_buffer, tmp_var);
      CONCAT_u32_u64_756_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_774_inst
    process(wp_buffer, wp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(wp_buffer, wp_buffer, tmp_var);
      CONCAT_u32_u64_774_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_776_call call_stmt_758_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_776_call_req_0;
      reqL_unguarded(0) <= call_stmt_758_call_req_0;
      call_stmt_776_call_ack_0 <= ackL_unguarded(1);
      call_stmt_758_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_776_call_req_1;
      reqR_unguarded(0) <= call_stmt_758_call_req_1;
      call_stmt_776_call_ack_1 <= ackR_unguarded(1);
      call_stmt_758_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_760_wire_constant & type_cast_762_wire_constant & CONCAT_u4_u8_768_wire_constant & ADD_u36_u36_771_wire & CONCAT_u32_u64_774_wire & type_cast_744_wire_constant & type_cast_746_wire_constant & CONCAT_u4_u8_752_wire_constant & q_base_address_buffer & CONCAT_u32_u64_756_wire;
      ignore_1_776 <= data_out(127 downto 64);
      ignore_758 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(31 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_3880_start: Boolean;
  signal transmitEngineDaemon_CP_3880_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_2196_branch_ack_0 : boolean;
  signal if_stmt_2196_branch_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_req_0 : boolean;
  signal phi_stmt_2216_req_0 : boolean;
  signal AND_u6_u6_2215_inst_req_0 : boolean;
  signal if_stmt_2196_branch_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_ack_0 : boolean;
  signal AND_u6_u6_2215_inst_ack_1 : boolean;
  signal AND_u6_u6_2215_inst_req_1 : boolean;
  signal AND_u6_u6_2215_inst_ack_0 : boolean;
  signal do_while_stmt_2204_branch_req_0 : boolean;
  signal phi_stmt_2216_req_1 : boolean;
  signal ncount_2290_2218_buf_ack_1 : boolean;
  signal ncount_2290_2218_buf_req_1 : boolean;
  signal ncount_2290_2218_buf_req_0 : boolean;
  signal ncount_2290_2218_buf_ack_0 : boolean;
  signal phi_stmt_2216_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_req_1 : boolean;
  signal call_stmt_2227_call_req_0 : boolean;
  signal call_stmt_2227_call_ack_0 : boolean;
  signal call_stmt_2227_call_req_1 : boolean;
  signal call_stmt_2227_call_ack_1 : boolean;
  signal call_stmt_2231_call_req_0 : boolean;
  signal call_stmt_2231_call_ack_0 : boolean;
  signal call_stmt_2231_call_req_1 : boolean;
  signal call_stmt_2231_call_ack_1 : boolean;
  signal NOT_u1_u1_2241_inst_req_0 : boolean;
  signal NOT_u1_u1_2241_inst_ack_0 : boolean;
  signal NOT_u1_u1_2241_inst_req_1 : boolean;
  signal NOT_u1_u1_2241_inst_ack_1 : boolean;
  signal W_pkt_pointer_2226_delayed_4_0_2251_inst_req_0 : boolean;
  signal W_pkt_pointer_2226_delayed_4_0_2251_inst_ack_0 : boolean;
  signal W_pkt_pointer_2226_delayed_4_0_2251_inst_req_1 : boolean;
  signal W_pkt_pointer_2226_delayed_4_0_2251_inst_ack_1 : boolean;
  signal call_stmt_2260_call_req_0 : boolean;
  signal call_stmt_2260_call_ack_0 : boolean;
  signal call_stmt_2260_call_req_1 : boolean;
  signal call_stmt_2260_call_ack_1 : boolean;
  signal W_count_2239_delayed_14_0_2264_inst_req_0 : boolean;
  signal W_count_2239_delayed_14_0_2264_inst_ack_0 : boolean;
  signal W_count_2239_delayed_14_0_2264_inst_req_1 : boolean;
  signal W_count_2239_delayed_14_0_2264_inst_ack_1 : boolean;
  signal call_stmt_2276_call_req_0 : boolean;
  signal call_stmt_2276_call_ack_0 : boolean;
  signal call_stmt_2276_call_req_1 : boolean;
  signal call_stmt_2276_call_ack_1 : boolean;
  signal ADD_u32_u32_2280_inst_req_0 : boolean;
  signal ADD_u32_u32_2280_inst_ack_0 : boolean;
  signal ADD_u32_u32_2280_inst_req_1 : boolean;
  signal ADD_u32_u32_2280_inst_ack_1 : boolean;
  signal W_count_2247_delayed_14_0_2282_inst_req_0 : boolean;
  signal W_count_2247_delayed_14_0_2282_inst_ack_0 : boolean;
  signal W_count_2247_delayed_14_0_2282_inst_req_1 : boolean;
  signal W_count_2247_delayed_14_0_2282_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_ack_1 : boolean;
  signal do_while_stmt_2204_branch_ack_0 : boolean;
  signal do_while_stmt_2204_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_3880_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3880_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3880_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3880_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_3880: Block -- control-path 
    signal transmitEngineDaemon_CP_3880_elements: BooleanArray(86 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_3880_elements(0) <= transmitEngineDaemon_CP_3880_start;
    transmitEngineDaemon_CP_3880_symbol <= transmitEngineDaemon_CP_3880_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_sample_start_
      -- CP-element group 0: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Sample/req
      -- CP-element group 0: 	 assign_stmt_2193/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Sample/$entry
      -- 
    req_3893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_sample_completed_
      -- CP-element group 1: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Update/$entry
      -- CP-element group 1: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_update_start_
      -- CP-element group 1: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Sample/ack
      -- CP-element group 1: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Update/req
      -- 
    ack_3894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(1)); -- 
    req_3898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	86 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_2194/$entry
      -- CP-element group 2: 	 assign_stmt_2193/$exit
      -- CP-element group 2: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2194/merge_stmt_2195__entry__
      -- CP-element group 2: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Update/ack
      -- CP-element group 2: 	 assign_stmt_2193/WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2194/branch_block_stmt_2194__entry__
      -- CP-element group 2: 	 branch_block_stmt_2194/merge_stmt_2195_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_2194/merge_stmt_2195__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_2194/merge_stmt_2195__entry___PhiReq/$exit
      -- 
    ack_3899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_2194/$exit
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_2194/branch_block_stmt_2194__exit__
      -- 
    transmitEngineDaemon_CP_3880_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	85 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	86 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_2194/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_2194/do_while_stmt_2204__exit__
      -- CP-element group 4: 	 branch_block_stmt_2194/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_2194/disable_loopback_PhiReq/$exit
      -- 
    transmitEngineDaemon_CP_3880_elements(4) <= transmitEngineDaemon_CP_3880_elements(85);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	86 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	86 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2194/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_2194/if_stmt_2196_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_2194/if_stmt_2196_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_2194/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_2194/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_3972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2196_branch_ack_1, ack => transmitEngineDaemon_CP_3880_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	86 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_2194/if_stmt_2196__exit__
      -- CP-element group 6: 	 branch_block_stmt_2194/do_while_stmt_2204__entry__
      -- CP-element group 6: 	 branch_block_stmt_2194/if_stmt_2196_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_2194/if_stmt_2196_else_link/else_choice_transition
      -- 
    else_choice_transition_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2196_branch_ack_0, ack => transmitEngineDaemon_CP_3880_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204__entry__
      -- CP-element group 7: 	 branch_block_stmt_2194/do_while_stmt_2204/$entry
      -- 
    transmitEngineDaemon_CP_3880_elements(7) <= transmitEngineDaemon_CP_3880_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	85 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204__exit__
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_back
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	83 
    -- CP-element group 10: 	84 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2194/do_while_stmt_2204/condition_done
      -- CP-element group 10: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_taken/$entry
      -- 
    transmitEngineDaemon_CP_3880_elements(10) <= transmitEngineDaemon_CP_3880_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	82 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_body_done
      -- 
    transmitEngineDaemon_CP_3880_elements(11) <= transmitEngineDaemon_CP_3880_elements(82);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/back_edge_to_loop_body
      -- 
    transmitEngineDaemon_CP_3880_elements(12) <= transmitEngineDaemon_CP_3880_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	31 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/first_time_through_loop_body
      -- 
    transmitEngineDaemon_CP_3880_elements(13) <= transmitEngineDaemon_CP_3880_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	25 
    -- CP-element group 14: 	26 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2206_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/$entry
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	81 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/condition_evaluated
      -- 
    condition_evaluated_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(15), ack => do_while_stmt_2204_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(81) & transmitEngineDaemon_CP_3880_elements(19);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	25 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_sample_start__ps
      -- CP-element group 16: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/aggregated_phi_sample_req
      -- 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(14) & transmitEngineDaemon_CP_3880_elements(25) & transmitEngineDaemon_CP_3880_elements(19);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	23 
    -- CP-element group 17: 	27 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	47 
    -- CP-element group 17: 	51 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	82 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	25 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2206_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/aggregated_phi_sample_ack
      -- 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(23) & transmitEngineDaemon_CP_3880_elements(27);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	26 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_update_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(20) & transmitEngineDaemon_CP_3880_elements(26);
      gj_transmitEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	28 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/aggregated_phi_update_ack
      -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(24) & transmitEngineDaemon_CP_3880_elements(28);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	44 
    -- CP-element group 20: 	79 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2206_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(14) & transmitEngineDaemon_CP_3880_elements(44) & transmitEngineDaemon_CP_3880_elements(79);
      gj_transmitEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Sample/$entry
      -- 
    rr_4009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(21), ack => AND_u6_u6_2215_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(16) & transmitEngineDaemon_CP_3880_elements(23);
      gj_transmitEngineDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_update_start_
      -- CP-element group 22: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Update/$entry
      -- 
    cr_4014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(22), ack => AND_u6_u6_2215_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(18) & transmitEngineDaemon_CP_3880_elements(24);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Sample/$exit
      -- 
    ra_4010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_2215_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	42 
    -- CP-element group 24: 	78 
    -- CP-element group 24: 	19 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2206_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/AND_u6_u6_2215_Update/$exit
      -- 
    ca_4015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_2215_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(24)); -- 
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	14 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	49 
    -- CP-element group 25: 	73 
    -- CP-element group 25: 	77 
    -- CP-element group 25: 	53 
    -- CP-element group 25: 	17 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_sample_start_
      -- 
    transmitEngineDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(14) & transmitEngineDaemon_CP_3880_elements(49) & transmitEngineDaemon_CP_3880_elements(73) & transmitEngineDaemon_CP_3880_elements(77) & transmitEngineDaemon_CP_3880_elements(53) & transmitEngineDaemon_CP_3880_elements(17);
      gj_transmitEngineDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	72 
    -- CP-element group 26: 	76 
    -- CP-element group 26: 	64 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	18 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(14) & transmitEngineDaemon_CP_3880_elements(72) & transmitEngineDaemon_CP_3880_elements(76) & transmitEngineDaemon_CP_3880_elements(64);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	17 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_sample_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28: 	62 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	19 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_update_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_loopback_trigger
      -- 
    transmitEngineDaemon_CP_3880_elements(29) <= transmitEngineDaemon_CP_3880_elements(12);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_loopback_sample_req
      -- CP-element group 30: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_loopback_sample_req_ps
      -- 
    phi_stmt_2216_loopback_sample_req_4025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2216_loopback_sample_req_4025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(30), ack => phi_stmt_2216_req_0); -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	13 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_entry_trigger
      -- 
    transmitEngineDaemon_CP_3880_elements(31) <= transmitEngineDaemon_CP_3880_elements(13);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_entry_sample_req
      -- CP-element group 32: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_entry_sample_req_ps
      -- 
    phi_stmt_2216_entry_sample_req_4028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2216_entry_sample_req_4028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(32), ack => phi_stmt_2216_req_1); -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_phi_mux_ack_ps
      -- CP-element group 33: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/phi_stmt_2216_phi_mux_ack
      -- 
    phi_stmt_2216_phi_mux_ack_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2216_ack_0, ack => transmitEngineDaemon_CP_3880_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Sample/req
      -- 
    req_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(34), ack => ncount_2290_2218_buf_req_0); -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_update_start_
      -- CP-element group 35: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Update/req
      -- 
    req_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(35), ack => ncount_2290_2218_buf_req_1); -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_sample_completed__ps
      -- 
    ack_4045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_2290_2218_buf_ack_0, ack => transmitEngineDaemon_CP_3880_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/R_ncount_2218_Update/$exit
      -- 
    ack_4050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_2290_2218_buf_ack_1, ack => transmitEngineDaemon_CP_3880_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_sample_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_update_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_update_completed__ps
      -- 
    transmitEngineDaemon_CP_3880_elements(40) <= transmitEngineDaemon_CP_3880_elements(41);
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	40 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/type_cast_2220_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3880_elements(39), ack => transmitEngineDaemon_CP_3880_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	24 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	69 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Sample/crr
      -- 
    crr_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(42), ack => call_stmt_2227_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(24) & transmitEngineDaemon_CP_3880_elements(44) & transmitEngineDaemon_CP_3880_elements(61) & transmitEngineDaemon_CP_3880_elements(69);
      gj_transmitEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	48 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	69 
    -- CP-element group 43: 	52 
    -- CP-element group 43: 	56 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_update_start_
      -- CP-element group 43: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Update/ccr
      -- 
    ccr_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(43), ack => call_stmt_2227_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(48) & transmitEngineDaemon_CP_3880_elements(61) & transmitEngineDaemon_CP_3880_elements(69) & transmitEngineDaemon_CP_3880_elements(52) & transmitEngineDaemon_CP_3880_elements(56);
      gj_transmitEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: 	20 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Sample/cra
      -- 
    cra_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2227_call_ack_0, ack => transmitEngineDaemon_CP_3880_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	50 
    -- CP-element group 45: 	54 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2227_Update/cca
      -- 
    cca_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2227_call_ack_1, ack => transmitEngineDaemon_CP_3880_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Sample/crr
      -- 
    crr_4081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(46), ack => call_stmt_2231_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(45) & transmitEngineDaemon_CP_3880_elements(48);
      gj_transmitEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	17 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	68 
    -- CP-element group 47: 	60 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_update_start_
      -- CP-element group 47: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Update/ccr
      -- 
    ccr_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(47), ack => call_stmt_2231_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(17) & transmitEngineDaemon_CP_3880_elements(68) & transmitEngineDaemon_CP_3880_elements(60);
      gj_transmitEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Sample/cra
      -- 
    cra_4082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2231_call_ack_0, ack => transmitEngineDaemon_CP_3880_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	66 
    -- CP-element group 49: 	58 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	25 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2231_Update/cca
      -- 
    cca_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2231_call_ack_1, ack => transmitEngineDaemon_CP_3880_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Sample/rr
      -- 
    rr_4095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(50), ack => NOT_u1_u1_2241_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(45) & transmitEngineDaemon_CP_3880_elements(52);
      gj_transmitEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	17 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	68 
    -- CP-element group 51: 	60 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_update_start_
      -- CP-element group 51: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Update/cr
      -- 
    cr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(51), ack => NOT_u1_u1_2241_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(17) & transmitEngineDaemon_CP_3880_elements(68) & transmitEngineDaemon_CP_3880_elements(60);
      gj_transmitEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	43 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Sample/ra
      -- 
    ra_4096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_2241_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	66 
    -- CP-element group 53: 	58 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	25 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/NOT_u1_u1_2241_Update/ca
      -- 
    ca_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_2241_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	45 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Sample/req
      -- 
    req_4109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(54), ack => W_pkt_pointer_2226_delayed_4_0_2251_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(45) & transmitEngineDaemon_CP_3880_elements(56);
      gj_transmitEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Update/req
      -- 
    req_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(55), ack => W_pkt_pointer_2226_delayed_4_0_2251_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3880_elements(60);
      gj_transmitEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Sample/ack
      -- 
    ack_4110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_2226_delayed_4_0_2251_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2253_Update/ack
      -- 
    ack_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_2226_delayed_4_0_2251_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Sample/crr
      -- 
    crr_4123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(58), ack => call_stmt_2260_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(49) & transmitEngineDaemon_CP_3880_elements(53) & transmitEngineDaemon_CP_3880_elements(57) & transmitEngineDaemon_CP_3880_elements(60);
      gj_transmitEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_update_start_
      -- CP-element group 59: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Update/ccr
      -- 
    ccr_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(59), ack => call_stmt_2260_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3880_elements(61);
      gj_transmitEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	47 
    -- CP-element group 60: 	51 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Sample/cra
      -- 
    cra_4124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2260_call_ack_0, ack => transmitEngineDaemon_CP_3880_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	82 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	42 
    -- CP-element group 61: 	43 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2260_Update/cca
      -- 
    cca_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2260_call_ack_1, ack => transmitEngineDaemon_CP_3880_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	28 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Sample/req
      -- 
    req_4137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(62), ack => W_count_2239_delayed_14_0_2264_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(28) & transmitEngineDaemon_CP_3880_elements(64);
      gj_transmitEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_update_start_
      -- CP-element group 63: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Update/req
      -- 
    req_4142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(63), ack => W_count_2239_delayed_14_0_2264_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3880_elements(68);
      gj_transmitEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	26 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Sample/ack
      -- 
    ack_4138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2239_delayed_14_0_2264_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2266_Update/ack
      -- 
    ack_4143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2239_delayed_14_0_2264_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	49 
    -- CP-element group 66: 	65 
    -- CP-element group 66: 	53 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Sample/crr
      -- 
    crr_4151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(66), ack => call_stmt_2276_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(49) & transmitEngineDaemon_CP_3880_elements(65) & transmitEngineDaemon_CP_3880_elements(53) & transmitEngineDaemon_CP_3880_elements(68);
      gj_transmitEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_update_start_
      -- CP-element group 67: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Update/ccr
      -- 
    ccr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(67), ack => call_stmt_2276_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3880_elements(69);
      gj_transmitEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	47 
    -- CP-element group 68: 	51 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Sample/cra
      -- 
    cra_4152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2276_call_ack_0, ack => transmitEngineDaemon_CP_3880_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	82 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	42 
    -- CP-element group 69: 	43 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/call_stmt_2276_Update/cca
      -- 
    cca_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2276_call_ack_1, ack => transmitEngineDaemon_CP_3880_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	28 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Sample/rr
      -- 
    rr_4165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(70), ack => ADD_u32_u32_2280_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(28) & transmitEngineDaemon_CP_3880_elements(72);
      gj_transmitEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_update_start_
      -- CP-element group 71: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Update/cr
      -- 
    cr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(71), ack => ADD_u32_u32_2280_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(17) & transmitEngineDaemon_CP_3880_elements(73);
      gj_transmitEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	26 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Sample/ra
      -- 
    ra_4166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2280_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	82 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	25 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/ADD_u32_u32_2280_Update/ca
      -- 
    ca_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2280_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Sample/req
      -- 
    req_4179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(74), ack => W_count_2247_delayed_14_0_2282_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(28) & transmitEngineDaemon_CP_3880_elements(76);
      gj_transmitEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Update/req
      -- 
    req_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(75), ack => W_count_2247_delayed_14_0_2282_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(17) & transmitEngineDaemon_CP_3880_elements(77);
      gj_transmitEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	26 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Sample/ack
      -- 
    ack_4180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2247_delayed_14_0_2282_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	25 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/assign_stmt_2284_Update/ack
      -- 
    ack_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2247_delayed_14_0_2282_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	24 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Sample/req
      -- 
    req_4193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(78), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(24) & transmitEngineDaemon_CP_3880_elements(80);
      gj_transmitEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	20 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Sample/ack
      -- CP-element group 79: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Update/req
      -- 
    ack_4194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_ack_0, ack => transmitEngineDaemon_CP_3880_elements(79)); -- 
    req_4198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(79), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_Update/ack
      -- 
    ack_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_ack_1, ack => transmitEngineDaemon_CP_3880_elements(80)); -- 
    -- CP-element group 81:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	15 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitEngineDaemon_CP_3880_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3880_elements(14), ack => transmitEngineDaemon_CP_3880_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  join  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	73 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	61 
    -- CP-element group 82: 	69 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	17 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	11 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2194/do_while_stmt_2204/do_while_stmt_2204_loop_body/$exit
      -- 
    transmitEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3880_elements(73) & transmitEngineDaemon_CP_3880_elements(77) & transmitEngineDaemon_CP_3880_elements(61) & transmitEngineDaemon_CP_3880_elements(69) & transmitEngineDaemon_CP_3880_elements(80) & transmitEngineDaemon_CP_3880_elements(17);
      gj_transmitEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	10 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_exit/$exit
      -- CP-element group 83: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_exit/ack
      -- 
    ack_4204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2204_branch_ack_0, ack => transmitEngineDaemon_CP_3880_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	10 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_taken/$exit
      -- CP-element group 84: 	 branch_block_stmt_2194/do_while_stmt_2204/loop_taken/ack
      -- 
    ack_4208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2204_branch_ack_1, ack => transmitEngineDaemon_CP_3880_elements(84)); -- 
    -- CP-element group 85:  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	4 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2194/do_while_stmt_2204/$exit
      -- 
    transmitEngineDaemon_CP_3880_elements(85) <= transmitEngineDaemon_CP_3880_elements(8);
    -- CP-element group 86:  merge  branch  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	2 
    -- CP-element group 86: 	4 
    -- CP-element group 86: 	5 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	5 
    -- CP-element group 86: 	6 
    -- CP-element group 86:  members (49) 
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196__entry__
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2194/merge_stmt_2195__exit__
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_else_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/NOT_u1_u1_2200_place
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Update/ack
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Update/req
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/BITSEL_u32_u1_2199/BITSEL_u32_u1_2199_inputs/RPIPE_CONTROL_REGISTER_2197/Sample/req
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_eval_test/NOT_u1_u1_2200/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/if_stmt_2196_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/merge_stmt_2195_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_2194/merge_stmt_2195_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_2194/merge_stmt_2195_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_2194/merge_stmt_2195_PhiAck/dummy
      -- 
    branch_req_3967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3880_elements(86), ack => if_stmt_2196_branch_req_0); -- 
    transmitEngineDaemon_CP_3880_elements(86) <= OrReduce(transmitEngineDaemon_CP_3880_elements(2) & transmitEngineDaemon_CP_3880_elements(4) & transmitEngineDaemon_CP_3880_elements(5));
    transmitEngineDaemon_do_while_stmt_2204_terminator_4209: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_2204_terminator_4209", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_3880_elements(11),loop_continue => transmitEngineDaemon_CP_3880_elements(84),loop_terminate => transmitEngineDaemon_CP_3880_elements(83),loop_back => transmitEngineDaemon_CP_3880_elements(9),loop_exit => transmitEngineDaemon_CP_3880_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_2216_phi_seq_4059_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitEngineDaemon_CP_3880_elements(29);
      transmitEngineDaemon_CP_3880_elements(34)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitEngineDaemon_CP_3880_elements(36);
      transmitEngineDaemon_CP_3880_elements(35)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitEngineDaemon_CP_3880_elements(37);
      transmitEngineDaemon_CP_3880_elements(30) <= phi_mux_reqs(0);
      triggers(1)  <= transmitEngineDaemon_CP_3880_elements(31);
      transmitEngineDaemon_CP_3880_elements(38)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitEngineDaemon_CP_3880_elements(38);
      transmitEngineDaemon_CP_3880_elements(39)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitEngineDaemon_CP_3880_elements(40);
      transmitEngineDaemon_CP_3880_elements(32) <= phi_mux_reqs(1);
      phi_stmt_2216_phi_seq_4059 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2216_phi_seq_4059") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitEngineDaemon_CP_3880_elements(16), 
          phi_sample_ack => transmitEngineDaemon_CP_3880_elements(27), 
          phi_update_req => transmitEngineDaemon_CP_3880_elements(18), 
          phi_update_ack => transmitEngineDaemon_CP_3880_elements(28), 
          phi_mux_ack => transmitEngineDaemon_CP_3880_elements(33), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3993_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_3880_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_3880_elements(13);
        entry_tmerge_3993 : transition_merge -- 
          generic map(name => " entry_tmerge_3993")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_3880_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_2246_2246_delayed_14_0_2281 : std_logic_vector(31 downto 0);
    signal ADD_u6_u6_2210_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_2215_wire : std_logic_vector(5 downto 0);
    signal BITSEL_u32_u1_2199_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2299_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2200_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2215_2215_delayed_4_0_2242 : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_2272_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_2197_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_2297_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_2257_wire : std_logic_vector(35 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_2208_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_2211_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_2213_wire : std_logic_vector(31 downto 0);
    signal count_2216 : std_logic_vector(31 downto 0);
    signal count_2239_delayed_14_0_2266 : std_logic_vector(31 downto 0);
    signal count_2247_delayed_14_0_2284 : std_logic_vector(31 downto 0);
    signal ignore_resp_2276 : std_logic_vector(31 downto 0);
    signal konst_2192_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2198_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2209_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2212_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2273_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2279_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2298_wire_constant : std_logic_vector(31 downto 0);
    signal ncount_2290 : std_logic_vector(31 downto 0);
    signal ncount_2290_2218_buffered : std_logic_vector(31 downto 0);
    signal pkt_pointer_2226_delayed_4_0_2253 : std_logic_vector(31 downto 0);
    signal pkt_pointer_2227 : std_logic_vector(31 downto 0);
    signal push_pointer_back_to_free_Q_2247 : std_logic_vector(0 downto 0);
    signal push_status_2260 : std_logic_vector(0 downto 0);
    signal transmitted_flag_2231 : std_logic_vector(0 downto 0);
    signal tx_flag_2227 : std_logic_vector(0 downto 0);
    signal tx_q_index_2206 : std_logic_vector(5 downto 0);
    signal type_cast_2214_wire : std_logic_vector(5 downto 0);
    signal type_cast_2220_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2256_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2269_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_2272_wire_constant <= "1111";
    konst_2192_wire_constant <= "000000";
    konst_2198_wire_constant <= "00000000000000000000000000000000";
    konst_2209_wire_constant <= "000001";
    konst_2212_wire_constant <= "00000000000000000000000000000001";
    konst_2273_wire_constant <= "010101";
    konst_2279_wire_constant <= "00000000000000000000000000000001";
    konst_2298_wire_constant <= "00000000000000000000000000000000";
    type_cast_2220_wire_constant <= "00000000000000000000000000000001";
    type_cast_2256_wire_constant <= "1";
    type_cast_2269_wire_constant <= "0";
    phi_stmt_2216: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ncount_2290_2218_buffered & type_cast_2220_wire_constant;
      req <= phi_stmt_2216_req_0 & phi_stmt_2216_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2216",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2216_ack_0,
          idata => idata,
          odata => count_2216,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2216
    -- flow-through select operator MUX_2289_inst
    ncount_2290 <= ADD_u32_u32_2246_2246_delayed_14_0_2281 when (push_pointer_back_to_free_Q_2247(0) /=  '0') else count_2247_delayed_14_0_2284;
    W_count_2239_delayed_14_0_2264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_2239_delayed_14_0_2264_inst_req_0;
      W_count_2239_delayed_14_0_2264_inst_ack_0<= wack(0);
      rreq(0) <= W_count_2239_delayed_14_0_2264_inst_req_1;
      W_count_2239_delayed_14_0_2264_inst_ack_1<= rack(0);
      W_count_2239_delayed_14_0_2264_inst : InterlockBuffer generic map ( -- 
        name => "W_count_2239_delayed_14_0_2264_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_2216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_2239_delayed_14_0_2266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_2247_delayed_14_0_2282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_2247_delayed_14_0_2282_inst_req_0;
      W_count_2247_delayed_14_0_2282_inst_ack_0<= wack(0);
      rreq(0) <= W_count_2247_delayed_14_0_2282_inst_req_1;
      W_count_2247_delayed_14_0_2282_inst_ack_1<= rack(0);
      W_count_2247_delayed_14_0_2282_inst : InterlockBuffer generic map ( -- 
        name => "W_count_2247_delayed_14_0_2282_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_2216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_2247_delayed_14_0_2284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_pointer_2226_delayed_4_0_2251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_pointer_2226_delayed_4_0_2251_inst_req_0;
      W_pkt_pointer_2226_delayed_4_0_2251_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_pointer_2226_delayed_4_0_2251_inst_req_1;
      W_pkt_pointer_2226_delayed_4_0_2251_inst_ack_1<= rack(0);
      W_pkt_pointer_2226_delayed_4_0_2251_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_pointer_2226_delayed_4_0_2251_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_pointer_2227,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_pointer_2226_delayed_4_0_2253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ncount_2290_2218_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_2290_2218_buf_req_0;
      ncount_2290_2218_buf_ack_0<= wack(0);
      rreq(0) <= ncount_2290_2218_buf_req_1;
      ncount_2290_2218_buf_ack_1<= rack(0);
      ncount_2290_2218_buf : InterlockBuffer generic map ( -- 
        name => "ncount_2290_2218_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_2290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_2290_2218_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2206
    process(AND_u6_u6_2215_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := AND_u6_u6_2215_wire(5 downto 0);
      tx_q_index_2206 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2214_inst
    process(SUB_u32_u32_2213_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_2213_wire(5 downto 0);
      type_cast_2214_wire <= tmp_var; -- 
    end process;
    do_while_stmt_2204_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_2299_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2204_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2204_branch_req_0,
          ack0 => do_while_stmt_2204_branch_ack_0,
          ack1 => do_while_stmt_2204_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2196_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2200_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2196_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2196_branch_req_0,
          ack0 => if_stmt_2196_branch_ack_0,
          ack1 => if_stmt_2196_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_2280_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= count_2216;
      ADD_u32_u32_2246_2246_delayed_14_0_2281 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2280_inst_req_0;
      ADD_u32_u32_2280_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2280_inst_req_1;
      ADD_u32_u32_2280_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u6_u6_2210_inst
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_2208_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_READ_TX_QUEUE_INDEX_2208_wire, konst_2209_wire_constant, tmp_var);
      ADD_u6_u6_2210_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2246_inst
    process(NOT_u1_u1_2215_2215_delayed_4_0_2242, transmitted_flag_2231) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_2215_2215_delayed_4_0_2242, transmitted_flag_2231, tmp_var);
      push_pointer_back_to_free_Q_2247 <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_2215_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_2210_wire & type_cast_2214_wire;
      AND_u6_u6_2215_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_2215_inst_req_0;
      AND_u6_u6_2215_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_2215_inst_req_1;
      AND_u6_u6_2215_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator BITSEL_u32_u1_2199_inst
    process(RPIPE_CONTROL_REGISTER_2197_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_2197_wire, konst_2198_wire_constant, tmp_var);
      BITSEL_u32_u1_2199_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_2299_inst
    process(RPIPE_CONTROL_REGISTER_2297_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_2297_wire, konst_2298_wire_constant, tmp_var);
      BITSEL_u32_u1_2299_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2200_inst
    process(BITSEL_u32_u1_2199_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_2199_wire, tmp_var);
      NOT_u1_u1_2200_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (7) : NOT_u1_u1_2241_inst 
    ApIntNot_group_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tx_flag_2227;
      NOT_u1_u1_2215_2215_delayed_4_0_2242 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_2241_inst_req_0;
      NOT_u1_u1_2241_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_2241_inst_req_1;
      NOT_u1_u1_2241_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_7_gI: SplitGuardInterface generic map(name => "ApIntNot_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u32_u32_2213_inst
    process(RPIPE_NUMBER_OF_SERVERS_2211_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_2211_wire, konst_2212_wire_constant, tmp_var);
      SUB_u32_u32_2213_wire <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_2197_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_2297_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_2257_wire <= FREE_Q;
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_2208_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_2211_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2191_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2192_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 6),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2293_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_2206;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2227_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2227_call_req_0;
      call_stmt_2227_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2227_call_req_1;
      call_stmt_2227_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_q_index_2206;
      pkt_pointer_2227 <= data_out(32 downto 1);
      tx_flag_2227 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(5 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(32 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2231_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2231_call_req_0;
      call_stmt_2231_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2231_call_req_1;
      call_stmt_2231_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not tx_flag_2227(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pkt_pointer_2227;
      transmitted_flag_2231 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(31 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2260_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2260_call_req_0;
      call_stmt_2260_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2260_call_req_1;
      call_stmt_2260_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_2247(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2256_wire_constant & RPIPE_FREE_Q_2257_wire & pkt_pointer_2226_delayed_4_0_2253;
      push_status_2260 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2276_call 
    AccessRegister_call_group_3: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2276_call_req_0;
      call_stmt_2276_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2276_call_req_1;
      call_stmt_2276_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_2247(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_3_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2269_wire_constant & NOT_u4_u4_2272_wire_constant & konst_2273_wire_constant & count_2239_delayed_14_0_2266;
      ignore_resp_2276 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    packet_pointer : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_call_acks : in   std_logic_vector(1 downto 0);
    accessMemory_call_data : out  std_logic_vector(219 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_return_acks : in   std_logic_vector(1 downto 0);
    accessMemory_return_data : in   std_logic_vector(127 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal packet_pointer_buffer :  std_logic_vector(31 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_3598_start: Boolean;
  signal transmitPacket_CP_3598_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_2079_call_req_0 : boolean;
  signal call_stmt_2079_call_ack_0 : boolean;
  signal call_stmt_2079_call_req_1 : boolean;
  signal call_stmt_2079_call_ack_1 : boolean;
  signal do_while_stmt_2092_branch_req_0 : boolean;
  signal phi_stmt_2094_req_1 : boolean;
  signal phi_stmt_2094_req_0 : boolean;
  signal phi_stmt_2094_ack_0 : boolean;
  signal SUB_u11_u11_2098_inst_req_0 : boolean;
  signal SUB_u11_u11_2098_inst_ack_0 : boolean;
  signal SUB_u11_u11_2098_inst_req_1 : boolean;
  signal SUB_u11_u11_2098_inst_ack_1 : boolean;
  signal ncount_down_2139_2099_buf_req_0 : boolean;
  signal ncount_down_2139_2099_buf_ack_0 : boolean;
  signal ncount_down_2139_2099_buf_req_1 : boolean;
  signal ncount_down_2139_2099_buf_ack_1 : boolean;
  signal phi_stmt_2100_req_1 : boolean;
  signal phi_stmt_2100_req_0 : boolean;
  signal phi_stmt_2100_ack_0 : boolean;
  signal ADD_u36_u36_2104_inst_req_0 : boolean;
  signal ADD_u36_u36_2104_inst_ack_0 : boolean;
  signal ADD_u36_u36_2104_inst_req_1 : boolean;
  signal ADD_u36_u36_2104_inst_ack_1 : boolean;
  signal nmem_addr_2144_2105_buf_req_0 : boolean;
  signal nmem_addr_2144_2105_buf_ack_0 : boolean;
  signal nmem_addr_2144_2105_buf_req_1 : boolean;
  signal nmem_addr_2144_2105_buf_ack_1 : boolean;
  signal call_stmt_2116_call_req_0 : boolean;
  signal call_stmt_2116_call_ack_0 : boolean;
  signal call_stmt_2116_call_req_1 : boolean;
  signal call_stmt_2116_call_ack_1 : boolean;
  signal CONCAT_u65_u73_2123_inst_req_0 : boolean;
  signal CONCAT_u65_u73_2123_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_2123_inst_req_1 : boolean;
  signal CONCAT_u65_u73_2123_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2117_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2117_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2117_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2117_inst_ack_1 : boolean;
  signal call_stmt_2134_call_req_0 : boolean;
  signal call_stmt_2134_call_ack_0 : boolean;
  signal call_stmt_2134_call_req_1 : boolean;
  signal call_stmt_2134_call_ack_1 : boolean;
  signal do_while_stmt_2092_branch_ack_0 : boolean;
  signal do_while_stmt_2092_branch_ack_1 : boolean;
  signal call_stmt_2169_call_req_0 : boolean;
  signal call_stmt_2169_call_ack_0 : boolean;
  signal call_stmt_2169_call_req_1 : boolean;
  signal call_stmt_2169_call_ack_1 : boolean;
  signal CONCAT_u65_u73_2178_inst_req_0 : boolean;
  signal CONCAT_u65_u73_2178_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_2178_inst_req_1 : boolean;
  signal CONCAT_u65_u73_2178_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2172_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2172_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2172_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2172_inst_ack_1 : boolean;
  signal EQ_u11_u1_2186_inst_req_0 : boolean;
  signal EQ_u11_u1_2186_inst_ack_0 : boolean;
  signal EQ_u11_u1_2186_inst_req_1 : boolean;
  signal EQ_u11_u1_2186_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_3598_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_3598_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_3598_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_3598_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_3598: Block -- control-path 
    signal transmitPacket_CP_3598_elements: BooleanArray(85 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_3598_elements(0) <= transmitPacket_CP_3598_start;
    transmitPacket_CP_3598_symbol <= transmitPacket_CP_3598_elements(85);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/$entry
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_sample_start_
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_update_start_
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Sample/crr
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Update/$entry
      -- CP-element group 0: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Update/ccr
      -- 
    ccr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(0), ack => call_stmt_2079_call_req_1); -- 
    crr_3611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(0), ack => call_stmt_2079_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_sample_completed_
      -- CP-element group 1: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Sample/cra
      -- 
    cra_3612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2079_call_ack_0, ack => transmitPacket_CP_3598_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_2066_to_assign_stmt_2087/$exit
      -- CP-element group 2: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_update_completed_
      -- CP-element group 2: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Update/$exit
      -- CP-element group 2: 	 assign_stmt_2066_to_assign_stmt_2087/call_stmt_2079_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_2091/$entry
      -- CP-element group 2: 	 branch_block_stmt_2091/branch_block_stmt_2091__entry__
      -- CP-element group 2: 	 branch_block_stmt_2091/do_while_stmt_2092__entry__
      -- 
    cca_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2079_call_ack_1, ack => transmitPacket_CP_3598_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	76 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	80 
    -- CP-element group 3: 	83 
    -- CP-element group 3: 	77 
    -- CP-element group 3: 	78 
    -- CP-element group 3: 	84 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_2091/do_while_stmt_2092__exit__
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187__entry__
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/$entry
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Update/cr
      -- 
    crr_3831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(3), ack => call_stmt_2169_call_req_0); -- 
    ccr_3836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(3), ack => call_stmt_2169_call_req_1); -- 
    cr_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(3), ack => CONCAT_u65_u73_2178_inst_req_1); -- 
    rr_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(3), ack => EQ_u11_u1_2186_inst_req_0); -- 
    cr_3878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(3), ack => EQ_u11_u1_2186_inst_req_1); -- 
    transmitPacket_CP_3598_elements(3) <= transmitPacket_CP_3598_elements(76);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_2091/do_while_stmt_2092/$entry
      -- CP-element group 4: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092__entry__
      -- 
    transmitPacket_CP_3598_elements(4) <= transmitPacket_CP_3598_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	76 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092__exit__
      -- 
    -- Element group transmitPacket_CP_3598_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_back
      -- 
    -- Element group transmitPacket_CP_3598_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	74 
    -- CP-element group 7: 	75 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_2091/do_while_stmt_2092/condition_done
      -- CP-element group 7: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_taken/$entry
      -- 
    transmitPacket_CP_3598_elements(7) <= transmitPacket_CP_3598_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	73 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_body_done
      -- 
    transmitPacket_CP_3598_elements(8) <= transmitPacket_CP_3598_elements(73);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	21 
    -- CP-element group 9: 	42 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/back_edge_to_loop_body
      -- 
    transmitPacket_CP_3598_elements(9) <= transmitPacket_CP_3598_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	44 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/first_time_through_loop_body
      -- 
    transmitPacket_CP_3598_elements(10) <= transmitPacket_CP_3598_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/loop_body_start
      -- 
    -- Element group transmitPacket_CP_3598_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	20 
    -- CP-element group 12: 	72 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/condition_evaluated
      -- 
    condition_evaluated_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(12), ack => do_while_stmt_2092_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(16) & transmitPacket_CP_3598_elements(20) & transmitPacket_CP_3598_elements(72);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	36 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_sample_start__ps
      -- 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(17) & transmitPacket_CP_3598_elements(36) & transmitPacket_CP_3598_elements(16);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	73 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	36 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_sample_completed_
      -- 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(19) & transmitPacket_CP_3598_elements(39);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	37 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	40 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/aggregated_phi_update_req
      -- CP-element group 15: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_update_start__ps
      -- 
    transmitPacket_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(18) & transmitPacket_CP_3598_elements(37);
      gj_transmitPacket_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	41 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/aggregated_phi_update_ack
      -- 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(20) & transmitPacket_CP_3598_elements(41);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_sample_start_
      -- 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(11) & transmitPacket_CP_3598_elements(14);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_update_start_
      -- 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(11) & transmitPacket_CP_3598_elements(20);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: 	12 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_loopback_trigger
      -- 
    transmitPacket_CP_3598_elements(21) <= transmitPacket_CP_3598_elements(9);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_loopback_sample_req_ps
      -- 
    phi_stmt_2094_loopback_sample_req_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2094_loopback_sample_req_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(22), ack => phi_stmt_2094_req_1); -- 
    -- Element group transmitPacket_CP_3598_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_entry_trigger
      -- 
    transmitPacket_CP_3598_elements(23) <= transmitPacket_CP_3598_elements(10);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_entry_sample_req_ps
      -- 
    phi_stmt_2094_entry_sample_req_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2094_entry_sample_req_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(24), ack => phi_stmt_2094_req_0); -- 
    -- Element group transmitPacket_CP_3598_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2094_phi_mux_ack_ps
      -- 
    phi_stmt_2094_phi_mux_ack_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2094_ack_0, ack => transmitPacket_CP_3598_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_update_start__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Sample/rr
      -- 
    rr_3675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(28), ack => SUB_u11_u11_2098_inst_req_0); -- 
    transmitPacket_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(26) & transmitPacket_CP_3598_elements(30);
      gj_transmitPacket_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_update_start_
      -- CP-element group 29: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Update/cr
      -- 
    cr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(29), ack => SUB_u11_u11_2098_inst_req_1); -- 
    transmitPacket_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(27) & transmitPacket_CP_3598_elements(31);
      gj_transmitPacket_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Sample/ra
      -- 
    ra_3676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u11_u11_2098_inst_ack_0, ack => transmitPacket_CP_3598_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/SUB_u11_u11_2098_Update/ca
      -- 
    ca_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u11_u11_2098_inst_ack_1, ack => transmitPacket_CP_3598_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Sample/req
      -- 
    req_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(32), ack => ncount_down_2139_2099_buf_req_0); -- 
    -- Element group transmitPacket_CP_3598_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_update_start_
      -- CP-element group 33: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Update/req
      -- 
    req_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(33), ack => ncount_down_2139_2099_buf_req_1); -- 
    -- Element group transmitPacket_CP_3598_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Sample/ack
      -- 
    ack_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_2139_2099_buf_ack_0, ack => transmitPacket_CP_3598_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_ncount_down_2099_Update/ack
      -- 
    ack_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_2139_2099_buf_ack_1, ack => transmitPacket_CP_3598_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	13 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_sample_start_
      -- 
    transmitPacket_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(11) & transmitPacket_CP_3598_elements(14);
      gj_transmitPacket_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	59 
    -- CP-element group 37: 	41 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	15 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_update_start_
      -- 
    transmitPacket_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(11) & transmitPacket_CP_3598_elements(70) & transmitPacket_CP_3598_elements(59) & transmitPacket_CP_3598_elements(41);
      gj_transmitPacket_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_sample_start__ps
      -- 
    transmitPacket_CP_3598_elements(38) <= transmitPacket_CP_3598_elements(13);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	15 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_update_start__ps
      -- 
    transmitPacket_CP_3598_elements(40) <= transmitPacket_CP_3598_elements(15);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	68 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	37 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	9 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_loopback_trigger
      -- 
    transmitPacket_CP_3598_elements(42) <= transmitPacket_CP_3598_elements(9);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_loopback_sample_req_ps
      -- 
    phi_stmt_2100_loopback_sample_req_3710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2100_loopback_sample_req_3710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(43), ack => phi_stmt_2100_req_1); -- 
    -- Element group transmitPacket_CP_3598_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	10 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_entry_trigger
      -- 
    transmitPacket_CP_3598_elements(44) <= transmitPacket_CP_3598_elements(10);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_entry_sample_req_ps
      -- 
    phi_stmt_2100_entry_sample_req_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2100_entry_sample_req_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(45), ack => phi_stmt_2100_req_0); -- 
    -- Element group transmitPacket_CP_3598_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/phi_stmt_2100_phi_mux_ack_ps
      -- 
    phi_stmt_2100_phi_mux_ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2100_ack_0, ack => transmitPacket_CP_3598_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_update_start__ps
      -- 
    -- Element group transmitPacket_CP_3598_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Sample/rr
      -- 
    rr_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(49), ack => ADD_u36_u36_2104_inst_req_0); -- 
    transmitPacket_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(47) & transmitPacket_CP_3598_elements(51);
      gj_transmitPacket_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_update_start_
      -- CP-element group 50: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Update/cr
      -- 
    cr_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(50), ack => ADD_u36_u36_2104_inst_req_1); -- 
    transmitPacket_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(48) & transmitPacket_CP_3598_elements(52);
      gj_transmitPacket_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Sample/ra
      -- 
    ra_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_2104_inst_ack_0, ack => transmitPacket_CP_3598_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/ADD_u36_u36_2104_Update/ca
      -- 
    ca_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_2104_inst_ack_1, ack => transmitPacket_CP_3598_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Sample/req
      -- 
    req_3747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(53), ack => nmem_addr_2144_2105_buf_req_0); -- 
    -- Element group transmitPacket_CP_3598_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_update_start__ps
      -- CP-element group 54: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_update_start_
      -- CP-element group 54: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Update/req
      -- 
    req_3752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(54), ack => nmem_addr_2144_2105_buf_req_1); -- 
    -- Element group transmitPacket_CP_3598_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Sample/ack
      -- 
    ack_3748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_2144_2105_buf_ack_0, ack => transmitPacket_CP_3598_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/R_nmem_addr_2105_Update/ack
      -- 
    ack_3753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_2144_2105_buf_ack_1, ack => transmitPacket_CP_3598_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Sample/crr
      -- 
    crr_3762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(57), ack => call_stmt_2116_call_req_0); -- 
    transmitPacket_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(41) & transmitPacket_CP_3598_elements(59);
      gj_transmitPacket_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	63 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_update_start_
      -- CP-element group 58: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Update/ccr
      -- 
    ccr_3767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(58), ack => call_stmt_2116_call_req_1); -- 
    transmitPacket_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(60) & transmitPacket_CP_3598_elements(63);
      gj_transmitPacket_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: 	37 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Sample/cra
      -- 
    cra_3763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2116_call_ack_0, ack => transmitPacket_CP_3598_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2116_Update/cca
      -- 
    cca_3768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2116_call_ack_1, ack => transmitPacket_CP_3598_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Sample/rr
      -- 
    rr_3776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(61), ack => CONCAT_u65_u73_2123_inst_req_0); -- 
    transmitPacket_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(60) & transmitPacket_CP_3598_elements(63);
      gj_transmitPacket_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	66 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Update/cr
      -- 
    cr_3781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(62), ack => CONCAT_u65_u73_2123_inst_req_1); -- 
    transmitPacket_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(64) & transmitPacket_CP_3598_elements(66);
      gj_transmitPacket_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	58 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Sample/ra
      -- 
    ra_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2123_inst_ack_0, ack => transmitPacket_CP_3598_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/CONCAT_u65_u73_2123_Update/ca
      -- 
    ca_3782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2123_inst_ack_1, ack => transmitPacket_CP_3598_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Sample/req
      -- 
    req_3790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(65), ack => WPIPE_nic_to_mac_transmit_pipe_2117_inst_req_0); -- 
    transmitPacket_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(64) & transmitPacket_CP_3598_elements(67);
      gj_transmitPacket_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	62 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Update/req
      -- 
    ack_3791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2117_inst_ack_0, ack => transmitPacket_CP_3598_elements(66)); -- 
    req_3795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(66), ack => WPIPE_nic_to_mac_transmit_pipe_2117_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	73 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/WPIPE_nic_to_mac_transmit_pipe_2117_Update/ack
      -- 
    ack_3796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2117_inst_ack_1, ack => transmitPacket_CP_3598_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	41 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Sample/crr
      -- 
    crr_3804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(68), ack => call_stmt_2134_call_req_0); -- 
    transmitPacket_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(41) & transmitPacket_CP_3598_elements(70);
      gj_transmitPacket_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Update/ccr
      -- 
    ccr_3809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(69), ack => call_stmt_2134_call_req_1); -- 
    transmitPacket_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitPacket_CP_3598_elements(71);
      gj_transmitPacket_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	37 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Sample/cra
      -- 
    cra_3805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2134_call_ack_0, ack => transmitPacket_CP_3598_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/call_stmt_2134_Update/cca
      -- 
    cca_3810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2134_call_ack_1, ack => transmitPacket_CP_3598_elements(71)); -- 
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	12 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitPacket_CP_3598_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => transmitPacket_CP_3598_elements(11), ack => transmitPacket_CP_3598_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	67 
    -- CP-element group 73: 	14 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	8 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2091/do_while_stmt_2092/do_while_stmt_2092_loop_body/$exit
      -- 
    transmitPacket_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(67) & transmitPacket_CP_3598_elements(14) & transmitPacket_CP_3598_elements(71);
      gj_transmitPacket_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	7 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_exit/$exit
      -- CP-element group 74: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_exit/ack
      -- 
    ack_3815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2092_branch_ack_0, ack => transmitPacket_CP_3598_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	7 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_taken/$exit
      -- CP-element group 75: 	 branch_block_stmt_2091/do_while_stmt_2092/loop_taken/ack
      -- 
    ack_3819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2092_branch_ack_1, ack => transmitPacket_CP_3598_elements(75)); -- 
    -- CP-element group 76:  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	5 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	3 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_2091/do_while_stmt_2092/$exit
      -- 
    transmitPacket_CP_3598_elements(76) <= transmitPacket_CP_3598_elements(5);
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	3 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Sample/cra
      -- 
    cra_3832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2169_call_ack_0, ack => transmitPacket_CP_3598_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	3 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/call_stmt_2169_Update/cca
      -- CP-element group 78: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Sample/rr
      -- 
    cca_3837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2169_call_ack_1, ack => transmitPacket_CP_3598_elements(78)); -- 
    rr_3845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(78), ack => CONCAT_u65_u73_2178_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Sample/ra
      -- 
    ra_3846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2178_inst_ack_0, ack => transmitPacket_CP_3598_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	3 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/CONCAT_u65_u73_2178_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Sample/req
      -- 
    ca_3851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2178_inst_ack_1, ack => transmitPacket_CP_3598_elements(80)); -- 
    req_3859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(80), ack => WPIPE_nic_to_mac_transmit_pipe_2172_inst_req_0); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_update_start_
      -- CP-element group 81: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Update/req
      -- 
    ack_3860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2172_inst_ack_0, ack => transmitPacket_CP_3598_elements(81)); -- 
    req_3864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3598_elements(81), ack => WPIPE_nic_to_mac_transmit_pipe_2172_inst_req_1); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/WPIPE_nic_to_mac_transmit_pipe_2172_Update/ack
      -- 
    ack_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2172_inst_ack_1, ack => transmitPacket_CP_3598_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	3 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Sample/ra
      -- 
    ra_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u11_u1_2186_inst_ack_0, ack => transmitPacket_CP_3598_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	3 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/EQ_u11_u1_2186_Update/ca
      -- 
    ca_3879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u11_u1_2186_inst_ack_1, ack => transmitPacket_CP_3598_elements(84)); -- 
    -- CP-element group 85:  join  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 $exit
      -- CP-element group 85: 	 branch_block_stmt_2091/$exit
      -- CP-element group 85: 	 branch_block_stmt_2091/branch_block_stmt_2091__exit__
      -- CP-element group 85: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187__exit__
      -- CP-element group 85: 	 branch_block_stmt_2091/call_stmt_2169_to_assign_stmt_2187/$exit
      -- 
    transmitPacket_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3598_elements(82) & transmitPacket_CP_3598_elements(84);
      gj_transmitPacket_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3598_elements(85), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_2092_terminator_3820: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_2092_terminator_3820", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_3598_elements(8),loop_continue => transmitPacket_CP_3598_elements(75),loop_terminate => transmitPacket_CP_3598_elements(74),loop_back => transmitPacket_CP_3598_elements(6),loop_exit => transmitPacket_CP_3598_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_2094_phi_seq_3700_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_3598_elements(23);
      transmitPacket_CP_3598_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_3598_elements(30);
      transmitPacket_CP_3598_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_3598_elements(31);
      transmitPacket_CP_3598_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_3598_elements(21);
      transmitPacket_CP_3598_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_3598_elements(34);
      transmitPacket_CP_3598_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_3598_elements(35);
      transmitPacket_CP_3598_elements(22) <= phi_mux_reqs(1);
      phi_stmt_2094_phi_seq_3700 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2094_phi_seq_3700") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_3598_elements(13), 
          phi_sample_ack => transmitPacket_CP_3598_elements(19), 
          phi_update_req => transmitPacket_CP_3598_elements(15), 
          phi_update_ack => transmitPacket_CP_3598_elements(20), 
          phi_mux_ack => transmitPacket_CP_3598_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2100_phi_seq_3754_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_3598_elements(44);
      transmitPacket_CP_3598_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_3598_elements(51);
      transmitPacket_CP_3598_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_3598_elements(52);
      transmitPacket_CP_3598_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_3598_elements(42);
      transmitPacket_CP_3598_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_3598_elements(55);
      transmitPacket_CP_3598_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_3598_elements(56);
      transmitPacket_CP_3598_elements(43) <= phi_mux_reqs(1);
      phi_stmt_2100_phi_seq_3754 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2100_phi_seq_3754") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_3598_elements(38), 
          phi_sample_ack => transmitPacket_CP_3598_elements(39), 
          phi_update_req => transmitPacket_CP_3598_elements(40), 
          phi_update_ack => transmitPacket_CP_3598_elements(41), 
          phi_mux_ack => transmitPacket_CP_3598_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3642_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_3598_elements(9);
        preds(1)  <= transmitPacket_CP_3598_elements(10);
        entry_tmerge_3642 : transition_merge -- 
          generic map(name => " entry_tmerge_3642")
          port map (preds => preds, symbol_out => transmitPacket_CP_3598_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_2104_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u1_u65_2121_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_2176_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u65_u73_2123_wire : std_logic_vector(72 downto 0);
    signal CONCAT_u65_u73_2178_wire : std_logic_vector(72 downto 0);
    signal NOT_u4_u4_2129_wire_constant : std_logic_vector(3 downto 0);
    signal R_FULL_BYTE_MASK_2074_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_2111_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_2122_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_2164_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u11_u11_2098_wire : std_logic_vector(10 downto 0);
    signal SUB_u36_u36_2184_wire : std_logic_vector(35 downto 0);
    signal control_data_2079 : std_logic_vector(63 downto 0);
    signal control_data_addr_2066 : std_logic_vector(35 downto 0);
    signal count_down_2094 : std_logic_vector(10 downto 0);
    signal data_2116 : std_logic_vector(63 downto 0);
    signal ignore_resp5_2134 : std_logic_vector(31 downto 0);
    signal konst_2097_wire_constant : std_logic_vector(10 downto 0);
    signal konst_2103_wire_constant : std_logic_vector(35 downto 0);
    signal konst_2130_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2137_wire_constant : std_logic_vector(10 downto 0);
    signal konst_2142_wire_constant : std_logic_vector(35 downto 0);
    signal konst_2153_wire_constant : std_logic_vector(10 downto 0);
    signal last_tkeep_2087 : std_logic_vector(7 downto 0);
    signal last_word_2169 : std_logic_vector(63 downto 0);
    signal mem_addr_2100 : std_logic_vector(35 downto 0);
    signal ncount_down_2139 : std_logic_vector(10 downto 0);
    signal ncount_down_2139_2099_buffered : std_logic_vector(10 downto 0);
    signal nmem_addr_2144 : std_logic_vector(35 downto 0);
    signal nmem_addr_2144_2105_buffered : std_logic_vector(35 downto 0);
    signal not_last_word_2155 : std_logic_vector(0 downto 0);
    signal packet_size_2083 : std_logic_vector(10 downto 0);
    signal slice_2132_wire : std_logic_vector(31 downto 0);
    signal type_cast_2071_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2073_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2077_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2108_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2110_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2114_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2119_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2126_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2161_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2163_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2167_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2174_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2185_wire : std_logic_vector(10 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_2129_wire_constant <= "1111";
    R_FULL_BYTE_MASK_2074_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_2111_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_2122_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_2164_wire_constant <= "11111111";
    konst_2097_wire_constant <= "00000010000";
    konst_2103_wire_constant <= "000000000000000000000000000000011000";
    konst_2130_wire_constant <= "110101";
    konst_2137_wire_constant <= "00000001000";
    konst_2142_wire_constant <= "000000000000000000000000000000001000";
    konst_2153_wire_constant <= "00000001000";
    type_cast_2071_wire_constant <= "0";
    type_cast_2073_wire_constant <= "1";
    type_cast_2077_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2108_wire_constant <= "0";
    type_cast_2110_wire_constant <= "1";
    type_cast_2114_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2119_wire_constant <= "0";
    type_cast_2126_wire_constant <= "0";
    type_cast_2161_wire_constant <= "0";
    type_cast_2163_wire_constant <= "1";
    type_cast_2167_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2174_wire_constant <= "1";
    phi_stmt_2094: Block -- phi operator 
      signal idata: std_logic_vector(21 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SUB_u11_u11_2098_wire & ncount_down_2139_2099_buffered;
      req <= phi_stmt_2094_req_0 & phi_stmt_2094_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2094",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 11) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2094_ack_0,
          idata => idata,
          odata => count_down_2094,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2094
    phi_stmt_2100: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_2104_wire & nmem_addr_2144_2105_buffered;
      req <= phi_stmt_2100_req_0 & phi_stmt_2100_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2100",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2100_ack_0,
          idata => idata,
          odata => mem_addr_2100,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2100
    -- flow-through slice operator slice_2082_inst
    packet_size_2083 <= control_data_2079(18 downto 8);
    -- flow-through slice operator slice_2086_inst
    last_tkeep_2087 <= control_data_2079(7 downto 0);
    -- flow-through slice operator slice_2132_inst
    slice_2132_wire <= mem_addr_2100(31 downto 0);
    ncount_down_2139_2099_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_2139_2099_buf_req_0;
      ncount_down_2139_2099_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_2139_2099_buf_req_1;
      ncount_down_2139_2099_buf_ack_1<= rack(0);
      ncount_down_2139_2099_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_2139_2099_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 11,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_2139,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_2139_2099_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmem_addr_2144_2105_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_2144_2105_buf_req_0;
      nmem_addr_2144_2105_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_2144_2105_buf_req_1;
      nmem_addr_2144_2105_buf_ack_1<= rack(0);
      nmem_addr_2144_2105_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_2144_2105_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_2144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_2144_2105_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2065_inst
    process(packet_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := packet_pointer_buffer(31 downto 0);
      control_data_addr_2066 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2185_inst
    process(SUB_u36_u36_2184_wire) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := SUB_u36_u36_2184_wire(10 downto 0);
      type_cast_2185_wire <= tmp_var; -- 
    end process;
    do_while_stmt_2092_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_2155;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2092_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2092_branch_req_0,
          ack0 => do_while_stmt_2092_branch_ack_0,
          ack1 => do_while_stmt_2092_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_2104_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= control_data_addr_2066;
      ADD_u36_u36_2104_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_2104_inst_req_0;
      ADD_u36_u36_2104_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_2104_inst_req_1;
      ADD_u36_u36_2104_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000011000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_2143_inst
    process(mem_addr_2100) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mem_addr_2100, konst_2142_wire_constant, tmp_var);
      nmem_addr_2144 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_2121_inst
    process(type_cast_2119_wire_constant, data_2116) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2119_wire_constant, data_2116, tmp_var);
      CONCAT_u1_u65_2121_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_2176_inst
    process(type_cast_2174_wire_constant, last_word_2169) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2174_wire_constant, last_word_2169, tmp_var);
      CONCAT_u1_u65_2176_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : CONCAT_u65_u73_2123_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_2121_wire;
      CONCAT_u65_u73_2123_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_2123_inst_req_0;
      CONCAT_u65_u73_2123_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_2123_inst_req_1;
      CONCAT_u65_u73_2123_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : CONCAT_u65_u73_2178_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_2176_wire & last_tkeep_2087;
      CONCAT_u65_u73_2178_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_2178_inst_req_0;
      CONCAT_u65_u73_2178_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_2178_inst_req_1;
      CONCAT_u65_u73_2178_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : EQ_u11_u1_2186_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_2083 & type_cast_2185_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u11_u1_2186_inst_req_0;
      EQ_u11_u1_2186_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u11_u1_2186_inst_req_1;
      EQ_u11_u1_2186_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : SUB_u11_u11_2098_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_2083;
      SUB_u11_u11_2098_wire <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u11_u11_2098_inst_req_0;
      SUB_u11_u11_2098_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u11_u11_2098_inst_req_1;
      SUB_u11_u11_2098_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000010000",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u11_u11_2138_inst
    process(count_down_2094) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_2094, konst_2137_wire_constant, tmp_var);
      ncount_down_2139 <= tmp_var; --
    end process;
    -- binary operator SUB_u36_u36_2184_inst
    process(nmem_addr_2144, control_data_addr_2066) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(nmem_addr_2144, control_data_addr_2066, tmp_var);
      SUB_u36_u36_2184_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u11_u1_2154_inst
    process(ncount_down_2139) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_2139, konst_2153_wire_constant, tmp_var);
      not_last_word_2155 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_2117_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2117_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_2117_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2117_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_2117_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_2123_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(1),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(1),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 73),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_to_mac_transmit_pipe_2172_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2172_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_2172_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2172_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_2172_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_2178_wire;
      nic_to_mac_transmit_pipe_write_1_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2169_call call_stmt_2079_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2169_call_req_0;
      reqL_unguarded(0) <= call_stmt_2079_call_req_0;
      call_stmt_2169_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2079_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2169_call_req_1;
      reqR_unguarded(0) <= call_stmt_2079_call_req_1;
      call_stmt_2169_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2079_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2161_wire_constant & type_cast_2163_wire_constant & R_FULL_BYTE_MASK_2164_wire_constant & nmem_addr_2144 & type_cast_2167_wire_constant & type_cast_2071_wire_constant & type_cast_2073_wire_constant & R_FULL_BYTE_MASK_2074_wire_constant & control_data_addr_2066 & type_cast_2077_wire_constant;
      last_word_2169 <= data_out(127 downto 64);
      control_data_2079 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(1),
          ackR => accessMemory_call_acks(1),
          dataR => accessMemory_call_data(219 downto 110),
          tagR => accessMemory_call_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(1), -- cross-over
          ackL => accessMemory_return_reqs(1), -- cross-over
          dataL => accessMemory_return_data(127 downto 64),
          tagL => accessMemory_return_tag(5 downto 3),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2116_call 
    accessMemory_call_group_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2116_call_req_0;
      call_stmt_2116_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2116_call_req_1;
      call_stmt_2116_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2108_wire_constant & type_cast_2110_wire_constant & R_FULL_BYTE_MASK_2111_wire_constant & mem_addr_2100 & type_cast_2114_wire_constant;
      data_2116 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2134_call 
    AccessRegister_call_group_2: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2134_call_req_0;
      call_stmt_2134_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2134_call_req_1;
      call_stmt_2134_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_2_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2126_wire_constant & NOT_u4_u4_2129_wire_constant & konst_2130_wire_constant & slice_2132_wire;
      ignore_resp5_2134 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity updateTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    updated_total_msgs : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity updateTotalMessages;
architecture updateTotalMessages_arch of updateTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal updated_total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal updated_total_msgs_update_enable: Boolean;
  -- output port buffer signals
  signal updateTotalMessages_CP_890_start: Boolean;
  signal updateTotalMessages_CP_890_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_796_call_req_0 : boolean;
  signal call_stmt_796_call_ack_1 : boolean;
  signal call_stmt_796_call_req_1 : boolean;
  signal call_stmt_796_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "updateTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= updated_total_msgs;
  updated_total_msgs_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  updateTotalMessages_CP_890_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "updateTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateTotalMessages_CP_890_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= updateTotalMessages_CP_890_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateTotalMessages_CP_890_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  updateTotalMessages_CP_890: Block -- control-path 
    signal updateTotalMessages_CP_890_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    updateTotalMessages_CP_890_elements(0) <= updateTotalMessages_CP_890_start;
    updateTotalMessages_CP_890_symbol <= updateTotalMessages_CP_890_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_796/$entry
      -- CP-element group 0: 	 call_stmt_796/call_stmt_796_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_796/call_stmt_796_sample_start_
      -- CP-element group 0: 	 call_stmt_796/call_stmt_796_Sample/crr
      -- CP-element group 0: 	 call_stmt_796/call_stmt_796_Sample/$entry
      -- CP-element group 0: 	 call_stmt_796/call_stmt_796_Update/ccr
      -- CP-element group 0: 	 call_stmt_796/call_stmt_796_Update/$entry
      -- 
    ccr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateTotalMessages_CP_890_elements(0), ack => call_stmt_796_call_req_1); -- 
    crr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateTotalMessages_CP_890_elements(0), ack => call_stmt_796_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_796/call_stmt_796_sample_completed_
      -- CP-element group 1: 	 call_stmt_796/call_stmt_796_Sample/$exit
      -- CP-element group 1: 	 call_stmt_796/call_stmt_796_Sample/cra
      -- 
    cra_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_796_call_ack_0, ack => updateTotalMessages_CP_890_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_796/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_796/call_stmt_796_update_completed_
      -- CP-element group 2: 	 call_stmt_796/call_stmt_796_Update/cca
      -- CP-element group 2: 	 call_stmt_796/call_stmt_796_Update/$exit
      -- 
    cca_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_796_call_ack_1, ack => updateTotalMessages_CP_890_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u32_u64_794_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_790_wire_constant : std_logic_vector(7 downto 0);
    signal rdata_796 : std_logic_vector(63 downto 0);
    signal type_cast_782_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_784_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_790_wire_constant <= "11110000";
    type_cast_782_wire_constant <= "0";
    type_cast_784_wire_constant <= "0";
    -- binary operator CONCAT_u32_u64_794_inst
    process(updated_total_msgs_buffer, updated_total_msgs_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(updated_total_msgs_buffer, updated_total_msgs_buffer, tmp_var);
      CONCAT_u32_u64_794_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_796_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_796_call_req_0;
      call_stmt_796_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_796_call_req_1;
      call_stmt_796_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_782_wire_constant & type_cast_784_wire_constant & CONCAT_u4_u8_790_wire_constant & q_base_address_buffer & CONCAT_u32_u64_794_wire;
      rdata_796 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end updateTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buffer_pointer : in  std_logic_vector(35 downto 0);
    packet_size : in  std_logic_vector(10 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 55)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(10 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_1412_start: Boolean;
  signal writeControlInformationToMem_CP_1412_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1191_call_req_0 : boolean;
  signal call_stmt_1191_call_ack_0 : boolean;
  signal call_stmt_1191_call_req_1 : boolean;
  signal call_stmt_1191_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 55) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(46 downto 36) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(46 downto 36);
  in_buffer_data_in(54 downto 47) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(54 downto 47);
  in_buffer_data_in(tag_length + 54 downto 55) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 54 downto 55);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_1412_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1412_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1412_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1412_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_1412: Block -- control-path 
    signal writeControlInformationToMem_CP_1412_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_1412_elements(0) <= writeControlInformationToMem_CP_1412_start;
    writeControlInformationToMem_CP_1412_symbol <= writeControlInformationToMem_CP_1412_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/$entry
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_sample_start_
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_update_start_
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Update/ccr
      -- 
    crr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_1412_elements(0), ack => call_stmt_1191_call_req_0); -- 
    ccr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_1412_elements(0), ack => call_stmt_1191_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Sample/cra
      -- 
    cra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1191_call_ack_0, ack => writeControlInformationToMem_CP_1412_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1182_to_call_stmt_1191/$exit
      -- CP-element group 2: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_update_completed_
      -- CP-element group 2: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1182_to_call_stmt_1191/call_stmt_1191_Update/cca
      -- 
    cca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1191_call_ack_1, ack => writeControlInformationToMem_CP_1412_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u11_u19_1180_wire : std_logic_vector(18 downto 0);
    signal R_FULL_BYTE_MASK_1187_wire_constant : std_logic_vector(7 downto 0);
    signal control_data_1182 : std_logic_vector(63 downto 0);
    signal ignore_return_1191 : std_logic_vector(63 downto 0);
    signal type_cast_1184_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1186_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1187_wire_constant <= "11111111";
    type_cast_1184_wire_constant <= "0";
    type_cast_1186_wire_constant <= "0";
    -- interlock type_cast_1181_inst
    process(CONCAT_u11_u19_1180_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 18 downto 0) := CONCAT_u11_u19_1180_wire(18 downto 0);
      control_data_1182 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u11_u19_1180_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(18 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u11_u19_1180_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1191_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1191_call_req_0;
      call_stmt_1191_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1191_call_req_1;
      call_stmt_1191_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1184_wire_constant & type_cast_1186_wire_constant & R_FULL_BYTE_MASK_1187_wire_constant & base_buffer_pointer_buffer & control_data_1182;
      ignore_return_1191 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf_pointer : in  std_logic_vector(35 downto 0);
    buf_position_out : out  std_logic_vector(35 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal buf_position_out_buffer :  std_logic_vector(35 downto 0);
  signal buf_position_out_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_1096_start: Boolean;
  signal writeEthernetHeaderToMem_CP_1096_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal nI_1078_1049_buf_req_0 : boolean;
  signal phi_stmt_1039_req_0 : boolean;
  signal nI_1078_1049_buf_ack_1 : boolean;
  signal do_while_stmt_1037_branch_req_0 : boolean;
  signal W_buf_position_out_1089_inst_req_1 : boolean;
  signal W_buf_position_out_1089_inst_ack_1 : boolean;
  signal RPIPE_nic_rx_to_header_1052_inst_ack_0 : boolean;
  signal phi_stmt_1045_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_1052_inst_req_0 : boolean;
  signal ADD_u36_u36_1043_inst_req_0 : boolean;
  signal phi_stmt_1045_req_1 : boolean;
  signal phi_stmt_1045_req_0 : boolean;
  signal ADD_u36_u36_1043_inst_ack_1 : boolean;
  signal phi_stmt_1039_req_1 : boolean;
  signal phi_stmt_1039_ack_0 : boolean;
  signal nI_1078_1049_buf_ack_0 : boolean;
  signal nI_1078_1049_buf_req_1 : boolean;
  signal RPIPE_nic_rx_to_header_1052_inst_ack_1 : boolean;
  signal ADD_u36_u36_1043_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_1052_inst_req_1 : boolean;
  signal nbuf_position_1083_1044_buf_ack_1 : boolean;
  signal nbuf_position_1083_1044_buf_req_1 : boolean;
  signal W_buf_position_out_1089_inst_ack_0 : boolean;
  signal W_buf_position_out_1089_inst_req_0 : boolean;
  signal nbuf_position_1083_1044_buf_ack_0 : boolean;
  signal do_while_stmt_1037_branch_ack_1 : boolean;
  signal nbuf_position_1083_1044_buf_req_0 : boolean;
  signal do_while_stmt_1037_branch_ack_0 : boolean;
  signal ADD_u36_u36_1043_inst_req_1 : boolean;
  signal call_stmt_1073_call_ack_1 : boolean;
  signal call_stmt_1073_call_req_1 : boolean;
  signal call_stmt_1073_call_ack_0 : boolean;
  signal call_stmt_1073_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_1096_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= buf_position_out_buffer;
  buf_position_out <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1096_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1096_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1096_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_1096: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_1096_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_1096_elements(0) <= writeEthernetHeaderToMem_CP_1096_start;
    writeEthernetHeaderToMem_CP_1096_symbol <= writeEthernetHeaderToMem_CP_1096_elements(68);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1036/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1036/do_while_stmt_1037__entry__
      -- CP-element group 0: 	 branch_block_stmt_1036/branch_block_stmt_1036__entry__
      -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	66 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	67 
    -- CP-element group 1: 	68 
    -- CP-element group 1:  members (10) 
      -- CP-element group 1: 	 assign_stmt_1091/assign_stmt_1091_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1091/assign_stmt_1091_Update/req
      -- CP-element group 1: 	 branch_block_stmt_1036/$exit
      -- CP-element group 1: 	 assign_stmt_1091/assign_stmt_1091_Sample/req
      -- CP-element group 1: 	 assign_stmt_1091/assign_stmt_1091_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_1091/assign_stmt_1091_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1036/do_while_stmt_1037__exit__
      -- CP-element group 1: 	 assign_stmt_1091/assign_stmt_1091_sample_start_
      -- CP-element group 1: 	 assign_stmt_1091/$entry
      -- CP-element group 1: 	 branch_block_stmt_1036/branch_block_stmt_1036__exit__
      -- 
    req_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(1), ack => W_buf_position_out_1089_inst_req_1); -- 
    req_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(1), ack => W_buf_position_out_1089_inst_req_0); -- 
    writeEthernetHeaderToMem_CP_1096_elements(1) <= writeEthernetHeaderToMem_CP_1096_elements(66);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1036/do_while_stmt_1037/$entry
      -- CP-element group 2: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037__entry__
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(2) <= writeEthernetHeaderToMem_CP_1096_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	66 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037__exit__
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_back
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	65 
    -- CP-element group 5: 	64 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1036/do_while_stmt_1037/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_exit/$entry
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(5) <= writeEthernetHeaderToMem_CP_1096_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	63 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_body_done
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(6) <= writeEthernetHeaderToMem_CP_1096_elements(63);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	40 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/back_edge_to_loop_body
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(7) <= writeEthernetHeaderToMem_CP_1096_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	42 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/first_time_through_loop_body
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(8) <= writeEthernetHeaderToMem_CP_1096_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	62 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1050_sample_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	62 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/condition_evaluated
      -- 
    condition_evaluated_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(10), ack => do_while_stmt_1037_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(14) & writeEthernetHeaderToMem_CP_1096_elements(62);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	54 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_sample_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(15) & writeEthernetHeaderToMem_CP_1096_elements(34) & writeEthernetHeaderToMem_CP_1096_elements(9) & writeEthernetHeaderToMem_CP_1096_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	56 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	63 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1050_sample_completed_
      -- 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(17) & writeEthernetHeaderToMem_CP_1096_elements(37) & writeEthernetHeaderToMem_CP_1096_elements(56);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	53 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	55 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_update_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(16) & writeEthernetHeaderToMem_CP_1096_elements(35) & writeEthernetHeaderToMem_CP_1096_elements(53);
      gj_writeEthernetHeaderToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	57 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/aggregated_phi_update_ack
      -- 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(18) & writeEthernetHeaderToMem_CP_1096_elements(39) & writeEthernetHeaderToMem_CP_1096_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(9) & writeEthernetHeaderToMem_CP_1096_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	60 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(9) & writeEthernetHeaderToMem_CP_1096_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	58 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(19) <= writeEthernetHeaderToMem_CP_1096_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_loopback_sample_req_ps
      -- 
    phi_stmt_1039_loopback_sample_req_1135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1039_loopback_sample_req_1135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(20), ack => phi_stmt_1039_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(21) <= writeEthernetHeaderToMem_CP_1096_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_entry_sample_req_ps
      -- 
    phi_stmt_1039_entry_sample_req_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1039_entry_sample_req_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(22), ack => phi_stmt_1039_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1039_phi_mux_ack
      -- 
    phi_stmt_1039_phi_mux_ack_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1039_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_sample_start_
      -- 
    rr_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(26), ack => ADD_u36_u36_1043_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(24) & writeEthernetHeaderToMem_CP_1096_elements(28);
      gj_writeEthernetHeaderToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Update/cr
      -- 
    cr_1159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(27), ack => ADD_u36_u36_1043_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(25) & writeEthernetHeaderToMem_CP_1096_elements(29);
      gj_writeEthernetHeaderToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Sample/ra
      -- 
    ra_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1043_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/ADD_u36_u36_1043_Update/$exit
      -- 
    ca_1160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1043_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Sample/req
      -- CP-element group 30: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Sample/$entry
      -- 
    req_1172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(30), ack => nbuf_position_1083_1044_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Update/req
      -- CP-element group 31: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_update_start_
      -- 
    req_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(31), ack => nbuf_position_1083_1044_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Sample/ack
      -- CP-element group 32: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_sample_completed_
      -- 
    ack_1173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1083_1044_buf_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Update/ack
      -- CP-element group 33: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nbuf_position_1044_update_completed_
      -- 
    ack_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1083_1044_buf_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(9) & writeEthernetHeaderToMem_CP_1096_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	39 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(9) & writeEthernetHeaderToMem_CP_1096_elements(39);
      gj_writeEthernetHeaderToMem_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_sample_start__ps
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(36) <= writeEthernetHeaderToMem_CP_1096_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_update_start__ps
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(38) <= writeEthernetHeaderToMem_CP_1096_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	35 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(40) <= writeEthernetHeaderToMem_CP_1096_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_loopback_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_loopback_sample_req
      -- 
    phi_stmt_1045_loopback_sample_req_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1045_loopback_sample_req_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(41), ack => phi_stmt_1045_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(42) <= writeEthernetHeaderToMem_CP_1096_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_entry_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_entry_sample_req
      -- 
    phi_stmt_1045_entry_sample_req_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1045_entry_sample_req_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(43), ack => phi_stmt_1045_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_phi_mux_ack_ps
      -- CP-element group 44: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1045_phi_mux_ack
      -- 
    phi_stmt_1045_phi_mux_ack_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1045_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(47) <= writeEthernetHeaderToMem_CP_1096_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/type_cast_1048_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1096_elements(46), ack => writeEthernetHeaderToMem_CP_1096_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_sample_start__ps
      -- 
    req_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(49), ack => nI_1078_1049_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Update/req
      -- CP-element group 50: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Update/$entry
      -- 
    req_1221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(50), ack => nI_1078_1049_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Sample/ack
      -- 
    ack_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_1078_1049_buf_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/R_nI_1049_Update/$exit
      -- 
    ack_1222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_1078_1049_buf_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	60 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1050_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(9) & writeEthernetHeaderToMem_CP_1096_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_sample_start_
      -- 
    rr_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(54), ack => RPIPE_nic_rx_to_header_1052_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(11) & writeEthernetHeaderToMem_CP_1096_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Update/cr
      -- 
    cr_1240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(55), ack => RPIPE_nic_rx_to_header_1052_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(56) & writeEthernetHeaderToMem_CP_1096_elements(13);
      gj_writeEthernetHeaderToMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_sample_completed_
      -- 
    ra_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_1052_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/RPIPE_nic_rx_to_header_1052_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/phi_stmt_1050_update_completed_
      -- 
    ca_1241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_1052_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Sample/crr
      -- CP-element group 58: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_sample_start_
      -- 
    crr_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(58), ack => call_stmt_1073_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(18) & writeEthernetHeaderToMem_CP_1096_elements(57) & writeEthernetHeaderToMem_CP_1096_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_update_start_
      -- 
    ccr_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1096_elements(59), ack => call_stmt_1073_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_1096_elements(61);
      gj_writeEthernetHeaderToMem_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	53 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Sample/cra
      -- CP-element group 60: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_sample_completed_
      -- 
    cra_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1073_call_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Update/cca
      -- CP-element group 61: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/call_stmt_1073_update_completed_
      -- 
    cca_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1073_call_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(61)); -- 
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	9 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	10 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1096_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1096_elements(9), ack => writeEthernetHeaderToMem_CP_1096_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	12 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	6 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1036/do_while_stmt_1037/do_while_stmt_1037_loop_body/$exit
      -- 
    writeEthernetHeaderToMem_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1096_elements(61) & writeEthernetHeaderToMem_CP_1096_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	5 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_exit/ack
      -- CP-element group 64: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_exit/$exit
      -- 
    ack_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1037_branch_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	5 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_taken/ack
      -- CP-element group 65: 	 branch_block_stmt_1036/do_while_stmt_1037/loop_taken/$exit
      -- 
    ack_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1037_branch_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(65)); -- 
    -- CP-element group 66:  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	1 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1036/do_while_stmt_1037/$exit
      -- 
    writeEthernetHeaderToMem_CP_1096_elements(66) <= writeEthernetHeaderToMem_CP_1096_elements(3);
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	1 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_1091/assign_stmt_1091_Sample/ack
      -- CP-element group 67: 	 assign_stmt_1091/assign_stmt_1091_Sample/$exit
      -- CP-element group 67: 	 assign_stmt_1091/assign_stmt_1091_sample_completed_
      -- 
    ack_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_buf_position_out_1089_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1096_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	1 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 assign_stmt_1091/assign_stmt_1091_Update/ack
      -- CP-element group 68: 	 assign_stmt_1091/assign_stmt_1091_Update/$exit
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 assign_stmt_1091/assign_stmt_1091_update_completed_
      -- CP-element group 68: 	 assign_stmt_1091/$exit
      -- 
    ack_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_buf_position_out_1089_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1096_elements(68)); -- 
    writeEthernetHeaderToMem_do_while_stmt_1037_terminator_1265: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_1037_terminator_1265", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_1096_elements(6),loop_continue => writeEthernetHeaderToMem_CP_1096_elements(65),loop_terminate => writeEthernetHeaderToMem_CP_1096_elements(64),loop_back => writeEthernetHeaderToMem_CP_1096_elements(4),loop_exit => writeEthernetHeaderToMem_CP_1096_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1039_phi_seq_1179_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_1096_elements(21);
      writeEthernetHeaderToMem_CP_1096_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_1096_elements(28);
      writeEthernetHeaderToMem_CP_1096_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_1096_elements(29);
      writeEthernetHeaderToMem_CP_1096_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_1096_elements(19);
      writeEthernetHeaderToMem_CP_1096_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_1096_elements(32);
      writeEthernetHeaderToMem_CP_1096_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_1096_elements(33);
      writeEthernetHeaderToMem_CP_1096_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1039_phi_seq_1179 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1039_phi_seq_1179") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_1096_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_1096_elements(17), 
          phi_update_req => writeEthernetHeaderToMem_CP_1096_elements(13), 
          phi_update_ack => writeEthernetHeaderToMem_CP_1096_elements(18), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_1096_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1045_phi_seq_1223_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_1096_elements(42);
      writeEthernetHeaderToMem_CP_1096_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_1096_elements(45);
      writeEthernetHeaderToMem_CP_1096_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_1096_elements(47);
      writeEthernetHeaderToMem_CP_1096_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_1096_elements(40);
      writeEthernetHeaderToMem_CP_1096_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_1096_elements(51);
      writeEthernetHeaderToMem_CP_1096_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_1096_elements(52);
      writeEthernetHeaderToMem_CP_1096_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1045_phi_seq_1223 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1045_phi_seq_1223") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_1096_elements(36), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_1096_elements(37), 
          phi_update_req => writeEthernetHeaderToMem_CP_1096_elements(38), 
          phi_update_ack => writeEthernetHeaderToMem_CP_1096_elements(39), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_1096_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1121_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_1096_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_1096_elements(8);
        entry_tmerge_1121 : transition_merge -- 
          generic map(name => " entry_tmerge_1121")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1096_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1043_wire : std_logic_vector(35 downto 0);
    signal I_1045 : std_logic_vector(3 downto 0);
    signal RPIPE_nic_rx_to_header_1052_wire : std_logic_vector(72 downto 0);
    signal ULE_u4_u1_1087_wire : std_logic_vector(0 downto 0);
    signal buf_position_1039 : std_logic_vector(35 downto 0);
    signal ethernet_header_1050 : std_logic_vector(72 downto 0);
    signal ignore_return_1073 : std_logic_vector(63 downto 0);
    signal konst_1042_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1076_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1081_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1086_wire_constant : std_logic_vector(3 downto 0);
    signal nI_1078 : std_logic_vector(3 downto 0);
    signal nI_1078_1049_buffered : std_logic_vector(3 downto 0);
    signal nbuf_position_1083 : std_logic_vector(35 downto 0);
    signal nbuf_position_1083_1044_buffered : std_logic_vector(35 downto 0);
    signal type_cast_1048_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1066_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1068_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_1060 : std_logic_vector(63 downto 0);
    signal wkeep_1064 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1042_wire_constant <= "000000000000000000000000000000001000";
    konst_1076_wire_constant <= "0001";
    konst_1081_wire_constant <= "000000000000000000000000000000001000";
    konst_1086_wire_constant <= "0001";
    type_cast_1048_wire_constant <= "0000";
    type_cast_1066_wire_constant <= "0";
    type_cast_1068_wire_constant <= "0";
    phi_stmt_1039: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1043_wire & nbuf_position_1083_1044_buffered;
      req <= phi_stmt_1039_req_0 & phi_stmt_1039_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1039",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1039_ack_0,
          idata => idata,
          odata => buf_position_1039,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1039
    phi_stmt_1045: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1048_wire_constant & nI_1078_1049_buffered;
      req <= phi_stmt_1045_req_0 & phi_stmt_1045_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1045",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1045_ack_0,
          idata => idata,
          odata => I_1045,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1045
    -- flow-through slice operator slice_1059_inst
    wdata_1060 <= ethernet_header_1050(71 downto 8);
    -- flow-through slice operator slice_1063_inst
    wkeep_1064 <= ethernet_header_1050(7 downto 0);
    W_buf_position_out_1089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_buf_position_out_1089_inst_req_0;
      W_buf_position_out_1089_inst_ack_0<= wack(0);
      rreq(0) <= W_buf_position_out_1089_inst_req_1;
      W_buf_position_out_1089_inst_ack_1<= rack(0);
      W_buf_position_out_1089_inst : InterlockBuffer generic map ( -- 
        name => "W_buf_position_out_1089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => buf_position_1039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => buf_position_out_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nI_1078_1049_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_1078_1049_buf_req_0;
      nI_1078_1049_buf_ack_0<= wack(0);
      rreq(0) <= nI_1078_1049_buf_req_1;
      nI_1078_1049_buf_ack_1<= rack(0);
      nI_1078_1049_buf : InterlockBuffer generic map ( -- 
        name => "nI_1078_1049_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_1078,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_1078_1049_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nbuf_position_1083_1044_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_1083_1044_buf_req_0;
      nbuf_position_1083_1044_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_1083_1044_buf_req_1;
      nbuf_position_1083_1044_buf_ack_1<= rack(0);
      nbuf_position_1083_1044_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_1083_1044_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_1083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_1083_1044_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1050
    process(RPIPE_nic_rx_to_header_1052_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_1052_wire(72 downto 0);
      ethernet_header_1050 <= tmp_var; -- 
    end process;
    do_while_stmt_1037_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULE_u4_u1_1087_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1037_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1037_branch_req_0,
          ack0 => do_while_stmt_1037_branch_ack_0,
          ack1 => do_while_stmt_1037_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1043_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_1043_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1043_inst_req_0;
      ADD_u36_u36_1043_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1043_inst_req_1;
      ADD_u36_u36_1043_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1082_inst
    process(buf_position_1039) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_1039, konst_1081_wire_constant, tmp_var);
      nbuf_position_1083 <= tmp_var; --
    end process;
    -- binary operator ADD_u4_u4_1077_inst
    process(I_1045) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_1045, konst_1076_wire_constant, tmp_var);
      nI_1078 <= tmp_var; --
    end process;
    -- binary operator ULE_u4_u1_1087_inst
    process(nI_1078) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(nI_1078, konst_1086_wire_constant, tmp_var);
      ULE_u4_u1_1087_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_1052_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_1052_inst_req_0;
      RPIPE_nic_rx_to_header_1052_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_1052_inst_req_1;
      RPIPE_nic_rx_to_header_1052_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_1052_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1073_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1073_call_req_0;
      call_stmt_1073_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1073_call_req_1;
      call_stmt_1073_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1066_wire_constant & type_cast_1068_wire_constant & wkeep_1064 & buf_position_1039 & wdata_1060;
      ignore_return_1073 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buf_pointer : in  std_logic_vector(35 downto 0);
    buf_pointer : in  std_logic_vector(35 downto 0);
    packet_size_32 : out  std_logic_vector(10 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 20)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_32_buffer :  std_logic_vector(10 downto 0);
  signal packet_size_32_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_1283_start: Boolean;
  signal writePayloadToMem_CP_1283_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u36_u36_1107_inst_req_0 : boolean;
  signal do_while_stmt_1101_branch_req_0 : boolean;
  signal phi_stmt_1103_ack_0 : boolean;
  signal ADD_u36_u36_1107_inst_ack_0 : boolean;
  signal ADD_u36_u36_1107_inst_ack_1 : boolean;
  signal ADD_u36_u36_1107_inst_req_1 : boolean;
  signal phi_stmt_1103_req_0 : boolean;
  signal phi_stmt_1103_req_1 : boolean;
  signal nbuf_position_1143_1108_buf_req_0 : boolean;
  signal nbuf_position_1143_1108_buf_ack_0 : boolean;
  signal nbuf_position_1143_1108_buf_req_1 : boolean;
  signal nbuf_position_1143_1108_buf_ack_1 : boolean;
  signal RPIPE_nic_rx_to_packet_1111_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1111_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1111_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_1111_inst_ack_1 : boolean;
  signal call_stmt_1138_call_req_0 : boolean;
  signal call_stmt_1138_call_ack_0 : boolean;
  signal call_stmt_1138_call_req_1 : boolean;
  signal call_stmt_1138_call_ack_1 : boolean;
  signal do_while_stmt_1101_branch_ack_0 : boolean;
  signal do_while_stmt_1101_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(71 downto 36) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 36);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_1283_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 20) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(10 downto 0) <= packet_size_32_buffer;
  packet_size_32 <= out_buffer_data_out(10 downto 0);
  out_buffer_data_in(11 downto 11) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(11 downto 11);
  out_buffer_data_in(19 downto 12) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(19 downto 12);
  out_buffer_data_in(tag_length + 19 downto 20) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 19 downto 20);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1283_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1283_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1283_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_1283: Block -- control-path 
    signal writePayloadToMem_CP_1283_elements: BooleanArray(47 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_1283_elements(0) <= writePayloadToMem_CP_1283_start;
    writePayloadToMem_CP_1283_symbol <= writePayloadToMem_CP_1283_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1100/do_while_stmt_1101__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1100/branch_block_stmt_1100__entry__
      -- CP-element group 0: 	 branch_block_stmt_1100/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	47 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1100/do_while_stmt_1101__exit__
      -- CP-element group 1: 	 branch_block_stmt_1100/branch_block_stmt_1100__exit__
      -- CP-element group 1: 	 branch_block_stmt_1100/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 assign_stmt_1156_to_assign_stmt_1171/$entry
      -- CP-element group 1: 	 assign_stmt_1156_to_assign_stmt_1171/$exit
      -- 
    writePayloadToMem_CP_1283_elements(1) <= writePayloadToMem_CP_1283_elements(47);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101__entry__
      -- CP-element group 2: 	 branch_block_stmt_1100/do_while_stmt_1101/$entry
      -- 
    writePayloadToMem_CP_1283_elements(2) <= writePayloadToMem_CP_1283_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	47 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101__exit__
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_back
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	45 
    -- CP-element group 5: 	46 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1100/do_while_stmt_1101/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_taken/$entry
      -- 
    writePayloadToMem_CP_1283_elements(5) <= writePayloadToMem_CP_1283_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	44 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_body_done
      -- 
    writePayloadToMem_CP_1283_elements(6) <= writePayloadToMem_CP_1283_elements(44);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/back_edge_to_loop_body
      -- 
    writePayloadToMem_CP_1283_elements(7) <= writePayloadToMem_CP_1283_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/first_time_through_loop_body
      -- 
    writePayloadToMem_CP_1283_elements(8) <= writePayloadToMem_CP_1283_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	43 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1109_sample_start_
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	43 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/condition_evaluated
      -- 
    condition_evaluated_1307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(10), ack => do_while_stmt_1101_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(43) & writePayloadToMem_CP_1283_elements(14);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	35 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_sample_start__ps
      -- 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(9) & writePayloadToMem_CP_1283_elements(15) & writePayloadToMem_CP_1283_elements(14);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	37 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	44 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1109_sample_completed_
      -- 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(17) & writePayloadToMem_CP_1283_elements(37);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	34 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_update_start__ps
      -- 
    writePayloadToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(16) & writePayloadToMem_CP_1283_elements(34);
      gj_writePayloadToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	38 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/aggregated_phi_update_ack
      -- 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(18) & writePayloadToMem_CP_1283_elements(38);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_sample_start_
      -- 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(9) & writePayloadToMem_CP_1283_elements(12);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_update_start_
      -- 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(9) & writePayloadToMem_CP_1283_elements(41);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_sample_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	39 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_update_completed_
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_loopback_trigger
      -- 
    writePayloadToMem_CP_1283_elements(19) <= writePayloadToMem_CP_1283_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_loopback_sample_req
      -- 
    phi_stmt_1103_loopback_sample_req_1322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1103_loopback_sample_req_1322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(20), ack => phi_stmt_1103_req_1); -- 
    -- Element group writePayloadToMem_CP_1283_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_entry_trigger
      -- 
    writePayloadToMem_CP_1283_elements(21) <= writePayloadToMem_CP_1283_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_entry_sample_req
      -- 
    phi_stmt_1103_entry_sample_req_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1103_entry_sample_req_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(22), ack => phi_stmt_1103_req_0); -- 
    -- Element group writePayloadToMem_CP_1283_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1103_phi_mux_ack_ps
      -- 
    phi_stmt_1103_phi_mux_ack_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1103_ack_0, ack => writePayloadToMem_CP_1283_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_sample_start_
      -- 
    rr_1341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(26), ack => ADD_u36_u36_1107_inst_req_0); -- 
    writePayloadToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(24) & writePayloadToMem_CP_1283_elements(28);
      gj_writePayloadToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Update/$entry
      -- 
    cr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(27), ack => ADD_u36_u36_1107_inst_req_1); -- 
    writePayloadToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(25) & writePayloadToMem_CP_1283_elements(29);
      gj_writePayloadToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_sample_completed_
      -- 
    ra_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1107_inst_ack_0, ack => writePayloadToMem_CP_1283_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/ADD_u36_u36_1107_Update/$exit
      -- 
    ca_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1107_inst_ack_1, ack => writePayloadToMem_CP_1283_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Sample/req
      -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(30), ack => nbuf_position_1143_1108_buf_req_0); -- 
    -- Element group writePayloadToMem_CP_1283_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Update/req
      -- 
    req_1364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(31), ack => nbuf_position_1143_1108_buf_req_1); -- 
    -- Element group writePayloadToMem_CP_1283_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Sample/ack
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1143_1108_buf_ack_0, ack => writePayloadToMem_CP_1283_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/R_nbuf_position_1108_Update/ack
      -- 
    ack_1365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1143_1108_buf_ack_1, ack => writePayloadToMem_CP_1283_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	41 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	13 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1109_update_start_
      -- 
    writePayloadToMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(9) & writePayloadToMem_CP_1283_elements(41);
      gj_writePayloadToMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Sample/rr
      -- 
    rr_1378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(35), ack => RPIPE_nic_rx_to_packet_1111_inst_req_0); -- 
    writePayloadToMem_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(11) & writePayloadToMem_CP_1283_elements(38);
      gj_writePayloadToMem_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: 	37 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_update_start_
      -- CP-element group 36: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Update/cr
      -- 
    cr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(36), ack => RPIPE_nic_rx_to_packet_1111_inst_req_1); -- 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(13) & writePayloadToMem_CP_1283_elements(37);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: 	36 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Sample/ra
      -- 
    ra_1379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1111_inst_ack_0, ack => writePayloadToMem_CP_1283_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	14 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	35 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/phi_stmt_1109_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/RPIPE_nic_rx_to_packet_1111_Update/ca
      -- 
    ca_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1111_inst_ack_1, ack => writePayloadToMem_CP_1283_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	18 
    -- CP-element group 39: 	38 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Sample/crr
      -- 
    crr_1392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(39), ack => call_stmt_1138_call_req_0); -- 
    writePayloadToMem_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(18) & writePayloadToMem_CP_1283_elements(38) & writePayloadToMem_CP_1283_elements(41);
      gj_writePayloadToMem_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Update/ccr
      -- 
    ccr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1283_elements(40), ack => call_stmt_1138_call_req_1); -- 
    writePayloadToMem_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_1283_elements(42);
      gj_writePayloadToMem_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	34 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Sample/cra
      -- 
    cra_1393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1138_call_ack_0, ack => writePayloadToMem_CP_1283_elements(41)); -- 
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/call_stmt_1138_Update/cca
      -- 
    cca_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1138_call_ack_1, ack => writePayloadToMem_CP_1283_elements(42)); -- 
    -- CP-element group 43:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	9 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	10 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writePayloadToMem_CP_1283_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_1283_elements(9), ack => writePayloadToMem_CP_1283_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: 	12 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	6 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1100/do_while_stmt_1101/do_while_stmt_1101_loop_body/$exit
      -- 
    writePayloadToMem_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1283_elements(42) & writePayloadToMem_CP_1283_elements(12);
      gj_writePayloadToMem_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	5 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_exit/$exit
      -- CP-element group 45: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_exit/ack
      -- 
    ack_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1101_branch_ack_0, ack => writePayloadToMem_CP_1283_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	5 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_taken/$exit
      -- CP-element group 46: 	 branch_block_stmt_1100/do_while_stmt_1101/loop_taken/ack
      -- 
    ack_1407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1101_branch_ack_1, ack => writePayloadToMem_CP_1283_elements(46)); -- 
    -- CP-element group 47:  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	3 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	1 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1100/do_while_stmt_1101/$exit
      -- 
    writePayloadToMem_CP_1283_elements(47) <= writePayloadToMem_CP_1283_elements(3);
    writePayloadToMem_do_while_stmt_1101_terminator_1408: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_1101_terminator_1408", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_1283_elements(6),loop_continue => writePayloadToMem_CP_1283_elements(46),loop_terminate => writePayloadToMem_CP_1283_elements(45),loop_back => writePayloadToMem_CP_1283_elements(4),loop_exit => writePayloadToMem_CP_1283_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1103_phi_seq_1366_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_1283_elements(21);
      writePayloadToMem_CP_1283_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_1283_elements(28);
      writePayloadToMem_CP_1283_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_1283_elements(29);
      writePayloadToMem_CP_1283_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_1283_elements(19);
      writePayloadToMem_CP_1283_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_1283_elements(32);
      writePayloadToMem_CP_1283_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_1283_elements(33);
      writePayloadToMem_CP_1283_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1103_phi_seq_1366 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1103_phi_seq_1366") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_1283_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_1283_elements(17), 
          phi_update_req => writePayloadToMem_CP_1283_elements(13), 
          phi_update_ack => writePayloadToMem_CP_1283_elements(18), 
          phi_mux_ack => writePayloadToMem_CP_1283_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1308_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_1283_elements(7);
        preds(1)  <= writePayloadToMem_CP_1283_elements(8);
        entry_tmerge_1308 : transition_merge -- 
          generic map(name => " entry_tmerge_1308")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_1283_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1107_wire : std_logic_vector(35 downto 0);
    signal EQ_u64_u1_1151_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1154_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1146_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_1111_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_1150_wire_constant : std_logic_vector(63 downto 0);
    signal SUB_u36_u36_1160_wire : std_logic_vector(35 downto 0);
    signal buf_position_1103 : std_logic_vector(35 downto 0);
    signal ignore_return_1138 : std_logic_vector(63 downto 0);
    signal konst_1106_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1141_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1153_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_1116 : std_logic_vector(0 downto 0);
    signal nbuf_position_1143 : std_logic_vector(35 downto 0);
    signal nbuf_position_1143_1108_buffered : std_logic_vector(35 downto 0);
    signal packet_size_11_1162 : std_logic_vector(10 downto 0);
    signal payload_data_1109 : std_logic_vector(72 downto 0);
    signal type_cast_1131_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_1120 : std_logic_vector(63 downto 0);
    signal wkeep_1124 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_1150_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    konst_1106_wire_constant <= "000000000000000000000000000000001000";
    konst_1141_wire_constant <= "000000000000000000000000000000001000";
    konst_1153_wire_constant <= "00000000";
    type_cast_1131_wire_constant <= "0";
    type_cast_1133_wire_constant <= "0";
    phi_stmt_1103: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1107_wire & nbuf_position_1143_1108_buffered;
      req <= phi_stmt_1103_req_0 & phi_stmt_1103_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1103",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1103_ack_0,
          idata => idata,
          odata => buf_position_1103,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1103
    -- flow-through slice operator slice_1115_inst
    last_bit_1116 <= payload_data_1109(72 downto 72);
    -- flow-through slice operator slice_1119_inst
    wdata_1120 <= payload_data_1109(71 downto 8);
    -- flow-through slice operator slice_1123_inst
    wkeep_1124 <= payload_data_1109(7 downto 0);
    -- interlock W_last_keep_1169_inst
    process(wkeep_1124) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_1124(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    -- interlock W_packet_size_32_1163_inst
    process(packet_size_11_1162) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := packet_size_11_1162(10 downto 0);
      packet_size_32_buffer <= tmp_var; -- 
    end process;
    nbuf_position_1143_1108_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_1143_1108_buf_req_0;
      nbuf_position_1143_1108_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_1143_1108_buf_req_1;
      nbuf_position_1143_1108_buf_ack_1<= rack(0);
      nbuf_position_1143_1108_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_1143_1108_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_1143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_1143_1108_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1109
    process(RPIPE_nic_rx_to_packet_1111_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_1111_wire(72 downto 0);
      payload_data_1109 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1161_inst
    process(SUB_u36_u36_1160_wire) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := SUB_u36_u36_1160_wire(10 downto 0);
      packet_size_11_1162 <= tmp_var; -- 
    end process;
    do_while_stmt_1101_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1146_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1101_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1101_branch_req_0,
          ack0 => do_while_stmt_1101_branch_ack_0,
          ack1 => do_while_stmt_1101_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1107_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_1107_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1107_inst_req_0;
      ADD_u36_u36_1107_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1107_inst_req_1;
      ADD_u36_u36_1107_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1142_inst
    process(buf_position_1103) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_1103, konst_1141_wire_constant, tmp_var);
      nbuf_position_1143 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1155_inst
    process(EQ_u64_u1_1151_wire, EQ_u8_u1_1154_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u64_u1_1151_wire, EQ_u8_u1_1154_wire, tmp_var);
      bad_packet_identifier_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1151_inst
    process(wdata_1120) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_1120, R_BAD_PACKET_DATA_1150_wire_constant, tmp_var);
      EQ_u64_u1_1151_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1154_inst
    process(wkeep_1124) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wkeep_1124, konst_1153_wire_constant, tmp_var);
      EQ_u8_u1_1154_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1146_inst
    process(last_bit_1116) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_1116, tmp_var);
      NOT_u1_u1_1146_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u36_u36_1160_inst
    process(buf_position_1103, base_buf_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(buf_position_1103, base_buf_pointer_buffer, tmp_var);
      SUB_u36_u36_1160_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_1111_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_1111_inst_req_0;
      RPIPE_nic_rx_to_packet_1111_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_1111_inst_req_1;
      RPIPE_nic_rx_to_packet_1111_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_1111_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1138_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1138_call_req_0;
      call_stmt_1138_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1138_call_req_1;
      call_stmt_1138_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1131_wire_constant & type_cast_1133_wire_constant & wkeep_1124 & buf_position_1103 & wdata_1120;
      ignore_return_1138 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    AFB_NIC_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
    AFB_NIC_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    enable_mac_pipe_read_data: out std_logic_vector(0 downto 0);
    enable_mac_pipe_read_req : in std_logic_vector(0 downto 0);
    enable_mac_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data: in std_logic_vector(72 downto 0);
    mac_to_nic_data_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(11 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(41 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(11 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(41 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(5 downto 0);
  -- declarations related to module AccessRegister
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module AccessRegister
  signal AccessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal AccessRegister_bmask :  std_logic_vector(3 downto 0);
  signal AccessRegister_register_index :  std_logic_vector(5 downto 0);
  signal AccessRegister_wdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_rdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_in_args    : std_logic_vector(42 downto 0);
  signal AccessRegister_out_args   : std_logic_vector(31 downto 0);
  signal AccessRegister_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal AccessRegister_tag_out   : std_logic_vector(4 downto 0);
  signal AccessRegister_start_req : std_logic;
  signal AccessRegister_start_ack : std_logic;
  signal AccessRegister_fin_req   : std_logic;
  signal AccessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module AccessRegister
  signal AccessRegister_call_reqs: std_logic_vector(6 downto 0);
  signal AccessRegister_call_acks: std_logic_vector(6 downto 0);
  signal AccessRegister_return_reqs: std_logic_vector(6 downto 0);
  signal AccessRegister_return_acks: std_logic_vector(6 downto 0);
  signal AccessRegister_call_data: std_logic_vector(300 downto 0);
  signal AccessRegister_call_tag: std_logic_vector(13 downto 0);
  signal AccessRegister_return_data: std_logic_vector(223 downto 0);
  signal AccessRegister_return_tag: std_logic_vector(13 downto 0);
  -- declarations related to module NicRegisterAccessDaemon
  component NicRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
      MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module NicRegisterAccessDaemon
  signal NicRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal NicRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal NicRegisterAccessDaemon_start_req : std_logic;
  signal NicRegisterAccessDaemon_start_ack : std_logic;
  signal NicRegisterAccessDaemon_fin_req   : std_logic;
  signal NicRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      FREE_Q : in std_logic_vector(35 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(35 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module SoftwareRegisterAccessDaemon
  component SoftwareRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      MAC_ENABLE : in std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      enable_mac_pipe_write_req : out  std_logic_vector(0 downto 0);
      enable_mac_pipe_write_ack : in   std_logic_vector(0 downto 0);
      enable_mac_pipe_write_data : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module SoftwareRegisterAccessDaemon
  signal SoftwareRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal SoftwareRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal SoftwareRegisterAccessDaemon_start_req : std_logic;
  signal SoftwareRegisterAccessDaemon_start_ack : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_req   : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module UpdateRegister
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module UpdateRegister
  signal UpdateRegister_bmask :  std_logic_vector(3 downto 0);
  signal UpdateRegister_rval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_wdata :  std_logic_vector(31 downto 0);
  signal UpdateRegister_index :  std_logic_vector(5 downto 0);
  signal UpdateRegister_wval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_in_args    : std_logic_vector(73 downto 0);
  signal UpdateRegister_out_args   : std_logic_vector(31 downto 0);
  signal UpdateRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal UpdateRegister_tag_out   : std_logic_vector(2 downto 0);
  signal UpdateRegister_start_req : std_logic;
  signal UpdateRegister_start_ack : std_logic;
  signal UpdateRegister_fin_req   : std_logic;
  signal UpdateRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module UpdateRegister
  signal UpdateRegister_call_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_data: std_logic_vector(147 downto 0);
  signal UpdateRegister_call_tag: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_data: std_logic_vector(63 downto 0);
  signal UpdateRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemory
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemory
  signal accessMemory_lock :  std_logic_vector(0 downto 0);
  signal accessMemory_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemory_bmask :  std_logic_vector(7 downto 0);
  signal accessMemory_addr :  std_logic_vector(35 downto 0);
  signal accessMemory_wdata :  std_logic_vector(63 downto 0);
  signal accessMemory_rdata :  std_logic_vector(63 downto 0);
  signal accessMemory_in_args    : std_logic_vector(109 downto 0);
  signal accessMemory_out_args   : std_logic_vector(63 downto 0);
  signal accessMemory_tag_in    : std_logic_vector(7 downto 0) := (others => '0');
  signal accessMemory_tag_out   : std_logic_vector(7 downto 0);
  signal accessMemory_start_req : std_logic;
  signal accessMemory_start_ack : std_logic;
  signal accessMemory_fin_req   : std_logic;
  signal accessMemory_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemory
  signal accessMemory_call_reqs: std_logic_vector(15 downto 0);
  signal accessMemory_call_acks: std_logic_vector(15 downto 0);
  signal accessMemory_return_reqs: std_logic_vector(15 downto 0);
  signal accessMemory_return_acks: std_logic_vector(15 downto 0);
  signal accessMemory_call_data: std_logic_vector(1759 downto 0);
  signal accessMemory_call_tag: std_logic_vector(47 downto 0);
  signal accessMemory_return_data: std_logic_vector(1023 downto 0);
  signal accessMemory_return_tag: std_logic_vector(47 downto 0);
  -- declarations related to module acquireLock
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireLock
  signal acquireLock_q_base_address :  std_logic_vector(35 downto 0);
  signal acquireLock_m_ok :  std_logic_vector(0 downto 0);
  signal acquireLock_in_args    : std_logic_vector(35 downto 0);
  signal acquireLock_out_args   : std_logic_vector(0 downto 0);
  signal acquireLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireLock_tag_out   : std_logic_vector(2 downto 0);
  signal acquireLock_start_req : std_logic;
  signal acquireLock_start_ack : std_logic;
  signal acquireLock_fin_req   : std_logic;
  signal acquireLock_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireLock
  signal acquireLock_call_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_call_acks: std_logic_vector(1 downto 0);
  signal acquireLock_return_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_return_acks: std_logic_vector(1 downto 0);
  signal acquireLock_call_data: std_logic_vector(71 downto 0);
  signal acquireLock_call_tag: std_logic_vector(1 downto 0);
  signal acquireLock_return_data: std_logic_vector(1 downto 0);
  signal acquireLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module delay_time
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueElement_read_index :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(31 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(67 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(31 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(67 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(31 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueueLength
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueLength
  signal getQueueLength_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueLength_Queue_Length :  std_logic_vector(31 downto 0);
  signal getQueueLength_in_args    : std_logic_vector(35 downto 0);
  signal getQueueLength_out_args   : std_logic_vector(31 downto 0);
  signal getQueueLength_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueueLength_tag_out   : std_logic_vector(2 downto 0);
  signal getQueueLength_start_req : std_logic;
  signal getQueueLength_start_ack : std_logic;
  signal getQueueLength_fin_req   : std_logic;
  signal getQueueLength_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueLength
  signal getQueueLength_call_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_call_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_return_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_return_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_call_data: std_logic_vector(71 downto 0);
  signal getQueueLength_call_tag: std_logic_vector(1 downto 0);
  signal getQueueLength_return_data: std_logic_vector(63 downto 0);
  signal getQueueLength_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(35 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(71 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTotalMessages
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTotalMessages
  signal getTotalMessages_q_base_address :  std_logic_vector(35 downto 0);
  signal getTotalMessages_total_msgs :  std_logic_vector(31 downto 0);
  signal getTotalMessages_in_args    : std_logic_vector(35 downto 0);
  signal getTotalMessages_out_args   : std_logic_vector(31 downto 0);
  signal getTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal getTotalMessages_start_req : std_logic;
  signal getTotalMessages_start_ack : std_logic;
  signal getTotalMessages_fin_req   : std_logic;
  signal getTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module getTotalMessages
  signal getTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_data: std_logic_vector(71 downto 0);
  signal getTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_data: std_logic_vector(63 downto 0);
  signal getTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_queue_index :  std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(31 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(54 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(35 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(35 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(1 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(1 downto 0);
      AccessRegister_call_data : out  std_logic_vector(85 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(1 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(1 downto 0);
      AccessRegister_return_data : in   std_logic_vector(63 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_lock :  std_logic_vector(0 downto 0);
  signal popFromQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(31 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(36 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(32 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(73 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(65 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(35 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(35 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_lock :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(31 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(68 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(206 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseLock
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseLock
  signal releaseLock_q_base_address :  std_logic_vector(35 downto 0);
  signal releaseLock_in_args    : std_logic_vector(35 downto 0);
  signal releaseLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseLock_tag_out   : std_logic_vector(2 downto 0);
  signal releaseLock_start_req : std_logic;
  signal releaseLock_start_ack : std_logic;
  signal releaseLock_fin_req   : std_logic;
  signal releaseLock_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseLock
  signal releaseLock_call_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_call_acks: std_logic_vector(1 downto 0);
  signal releaseLock_return_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_return_acks: std_logic_vector(1 downto 0);
  signal releaseLock_call_data: std_logic_vector(71 downto 0);
  signal releaseLock_call_tag: std_logic_vector(1 downto 0);
  signal releaseLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueueElement_write_index :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(31 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(99 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(99 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(99 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(199 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(31 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_packet_pointer :  std_logic_vector(31 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(31 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(31 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module updateTotalMessages
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module updateTotalMessages
  signal updateTotalMessages_q_base_address :  std_logic_vector(35 downto 0);
  signal updateTotalMessages_updated_total_msgs :  std_logic_vector(31 downto 0);
  signal updateTotalMessages_in_args    : std_logic_vector(67 downto 0);
  signal updateTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal updateTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal updateTotalMessages_start_req : std_logic;
  signal updateTotalMessages_start_ack : std_logic;
  signal updateTotalMessages_fin_req   : std_logic;
  signal updateTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module updateTotalMessages
  signal updateTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal updateTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal updateTotalMessages_call_data: std_logic_vector(135 downto 0);
  signal updateTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(10 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(35 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(10 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(54 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(54 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position_out : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_buf_position_out :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(10 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_packet_size_32 :  std_logic_vector(10 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(71 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(19 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(71 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(19 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe CONTROL_REGISTER
  signal CONTROL_REGISTER_pipe_write_data: std_logic_vector(31 downto 0);
  signal CONTROL_REGISTER_pipe_write_req: std_logic_vector(0 downto 0);
  signal CONTROL_REGISTER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe CONTROL_REGISTER
  signal CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe FREE_Q
  signal FREE_Q_pipe_write_data: std_logic_vector(35 downto 0);
  signal FREE_Q_pipe_write_req: std_logic_vector(0 downto 0);
  signal FREE_Q_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe FREE_Q
  signal FREE_Q: std_logic_vector(35 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe MAC_ENABLE
  signal MAC_ENABLE_pipe_write_data: std_logic_vector(0 downto 0);
  signal MAC_ENABLE_pipe_write_req: std_logic_vector(0 downto 0);
  signal MAC_ENABLE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe MAC_ENABLE
  signal MAC_ENABLE: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(31 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(0 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe enable_mac
  signal enable_mac_pipe_write_data: std_logic_vector(0 downto 0);
  signal enable_mac_pipe_write_req: std_logic_vector(0 downto 0);
  signal enable_mac_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(145 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module AccessRegister
  AccessRegister_rwbar <= AccessRegister_in_args(42 downto 42);
  AccessRegister_bmask <= AccessRegister_in_args(41 downto 38);
  AccessRegister_register_index <= AccessRegister_in_args(37 downto 32);
  AccessRegister_wdata <= AccessRegister_in_args(31 downto 0);
  AccessRegister_out_args <= AccessRegister_rdata ;
  -- call arbiter for module AccessRegister
  AccessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 7,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => AccessRegister_call_reqs,
      call_acks => AccessRegister_call_acks,
      return_reqs => AccessRegister_return_reqs,
      return_acks => AccessRegister_return_acks,
      call_data  => AccessRegister_call_data,
      call_tag  => AccessRegister_call_tag,
      return_tag  => AccessRegister_return_tag,
      call_mtag => AccessRegister_tag_in,
      return_mtag => AccessRegister_tag_out,
      return_data =>AccessRegister_return_data,
      call_mreq => AccessRegister_start_req,
      call_mack => AccessRegister_start_ack,
      return_mreq => AccessRegister_fin_req,
      return_mack => AccessRegister_fin_ack,
      call_mdata => AccessRegister_in_args,
      return_mdata => AccessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  AccessRegister_instance:AccessRegister-- 
    generic map(tag_length => 5)
    port map(-- 
      rwbar => AccessRegister_rwbar,
      bmask => AccessRegister_bmask,
      register_index => AccessRegister_register_index,
      wdata => AccessRegister_wdata,
      rdata => AccessRegister_rdata,
      start_req => AccessRegister_start_req,
      start_ack => AccessRegister_start_ack,
      fin_req => AccessRegister_fin_req,
      fin_ack => AccessRegister_fin_ack,
      clk => clk,
      reset => reset,
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
      tag_in => AccessRegister_tag_in,
      tag_out => AccessRegister_tag_out-- 
    ); -- 
  -- module NicRegisterAccessDaemon
  NicRegisterAccessDaemon_instance:NicRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => NicRegisterAccessDaemon_start_req,
      start_ack => NicRegisterAccessDaemon_start_ack,
      fin_req => NicRegisterAccessDaemon_fin_req,
      fin_ack => NicRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(11 downto 6),
      memory_space_0_lr_tag => memory_space_0_lr_tag(41 downto 21),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(5 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(20 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
      MAC_ENABLE_pipe_write_req => MAC_ENABLE_pipe_write_req(0 downto 0),
      MAC_ENABLE_pipe_write_ack => MAC_ENABLE_pipe_write_ack(0 downto 0),
      MAC_ENABLE_pipe_write_data => MAC_ENABLE_pipe_write_data(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(1 downto 1),
      UpdateRegister_call_acks => UpdateRegister_call_acks(1 downto 1),
      UpdateRegister_call_data => UpdateRegister_call_data(147 downto 74),
      UpdateRegister_call_tag => UpdateRegister_call_tag(1 downto 1),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(1 downto 1),
      UpdateRegister_return_acks => UpdateRegister_return_acks(1 downto 1),
      UpdateRegister_return_data => UpdateRegister_return_data(63 downto 32),
      UpdateRegister_return_tag => UpdateRegister_return_tag(1 downto 1),
      tag_in => NicRegisterAccessDaemon_tag_in,
      tag_out => NicRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  NicRegisterAccessDaemon_tag_in <= (others => '0');
  NicRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => NicRegisterAccessDaemon_start_req, start_ack => NicRegisterAccessDaemon_start_ack,  fin_req => NicRegisterAccessDaemon_fin_req,  fin_ack => NicRegisterAccessDaemon_fin_ack);
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      FREE_Q => FREE_Q,
      CONTROL_REGISTER => CONTROL_REGISTER,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(5 downto 5),
      AccessRegister_call_acks => AccessRegister_call_acks(5 downto 5),
      AccessRegister_call_data => AccessRegister_call_data(257 downto 215),
      AccessRegister_call_tag => AccessRegister_call_tag(11 downto 10),
      AccessRegister_return_reqs => AccessRegister_return_reqs(5 downto 5),
      AccessRegister_return_acks => AccessRegister_return_acks(5 downto 5),
      AccessRegister_return_data => AccessRegister_return_data(191 downto 160),
      AccessRegister_return_tag => AccessRegister_return_tag(11 downto 10),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(73 downto 37),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(65 downto 33),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(35 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(137 downto 69),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(35 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module SoftwareRegisterAccessDaemon
  SoftwareRegisterAccessDaemon_instance:SoftwareRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => SoftwareRegisterAccessDaemon_start_req,
      start_ack => SoftwareRegisterAccessDaemon_start_ack,
      fin_req => SoftwareRegisterAccessDaemon_fin_req,
      fin_ack => SoftwareRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(5 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(20 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      MAC_ENABLE => MAC_ENABLE,
      FREE_Q_pipe_write_req => FREE_Q_pipe_write_req(0 downto 0),
      FREE_Q_pipe_write_ack => FREE_Q_pipe_write_ack(0 downto 0),
      FREE_Q_pipe_write_data => FREE_Q_pipe_write_data(35 downto 0),
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      CONTROL_REGISTER_pipe_write_req => CONTROL_REGISTER_pipe_write_req(0 downto 0),
      CONTROL_REGISTER_pipe_write_ack => CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      CONTROL_REGISTER_pipe_write_data => CONTROL_REGISTER_pipe_write_data(31 downto 0),
      NUMBER_OF_SERVERS_pipe_write_req => NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_ack => NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_data => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      enable_mac_pipe_write_req => enable_mac_pipe_write_req(0 downto 0),
      enable_mac_pipe_write_ack => enable_mac_pipe_write_ack(0 downto 0),
      enable_mac_pipe_write_data => enable_mac_pipe_write_data(0 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(0 downto 0),
      UpdateRegister_call_acks => UpdateRegister_call_acks(0 downto 0),
      UpdateRegister_call_data => UpdateRegister_call_data(73 downto 0),
      UpdateRegister_call_tag => UpdateRegister_call_tag(0 downto 0),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(0 downto 0),
      UpdateRegister_return_acks => UpdateRegister_return_acks(0 downto 0),
      UpdateRegister_return_data => UpdateRegister_return_data(31 downto 0),
      UpdateRegister_return_tag => UpdateRegister_return_tag(0 downto 0),
      tag_in => SoftwareRegisterAccessDaemon_tag_in,
      tag_out => SoftwareRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  SoftwareRegisterAccessDaemon_tag_in <= (others => '0');
  SoftwareRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => SoftwareRegisterAccessDaemon_start_req, start_ack => SoftwareRegisterAccessDaemon_start_ack,  fin_req => SoftwareRegisterAccessDaemon_fin_req,  fin_ack => SoftwareRegisterAccessDaemon_fin_ack);
  -- module UpdateRegister
  UpdateRegister_bmask <= UpdateRegister_in_args(73 downto 70);
  UpdateRegister_rval <= UpdateRegister_in_args(69 downto 38);
  UpdateRegister_wdata <= UpdateRegister_in_args(37 downto 6);
  UpdateRegister_index <= UpdateRegister_in_args(5 downto 0);
  UpdateRegister_out_args <= UpdateRegister_wval ;
  -- call arbiter for module UpdateRegister
  UpdateRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 74,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => UpdateRegister_call_reqs,
      call_acks => UpdateRegister_call_acks,
      return_reqs => UpdateRegister_return_reqs,
      return_acks => UpdateRegister_return_acks,
      call_data  => UpdateRegister_call_data,
      call_tag  => UpdateRegister_call_tag,
      return_tag  => UpdateRegister_return_tag,
      call_mtag => UpdateRegister_tag_in,
      return_mtag => UpdateRegister_tag_out,
      return_data =>UpdateRegister_return_data,
      call_mreq => UpdateRegister_start_req,
      call_mack => UpdateRegister_start_ack,
      return_mreq => UpdateRegister_fin_req,
      return_mack => UpdateRegister_fin_ack,
      call_mdata => UpdateRegister_in_args,
      return_mdata => UpdateRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  UpdateRegister_instance:UpdateRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      bmask => UpdateRegister_bmask,
      rval => UpdateRegister_rval,
      wdata => UpdateRegister_wdata,
      index => UpdateRegister_index,
      wval => UpdateRegister_wval,
      start_req => UpdateRegister_start_req,
      start_ack => UpdateRegister_start_ack,
      fin_req => UpdateRegister_fin_req,
      fin_ack => UpdateRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(11 downto 6),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 32),
      memory_space_0_sr_tag => memory_space_0_sr_tag(41 downto 21),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(5 downto 3),
      tag_in => UpdateRegister_tag_in,
      tag_out => UpdateRegister_tag_out-- 
    ); -- 
  -- module accessMemory
  accessMemory_lock <= accessMemory_in_args(109 downto 109);
  accessMemory_rwbar <= accessMemory_in_args(108 downto 108);
  accessMemory_bmask <= accessMemory_in_args(107 downto 100);
  accessMemory_addr <= accessMemory_in_args(99 downto 64);
  accessMemory_wdata <= accessMemory_in_args(63 downto 0);
  accessMemory_out_args <= accessMemory_rdata ;
  -- call arbiter for module accessMemory
  accessMemory_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 16,
      call_data_width => 110,
      return_data_width => 64,
      callee_tag_length => 5,
      caller_tag_length => 3--
    )
    port map(-- 
      call_reqs => accessMemory_call_reqs,
      call_acks => accessMemory_call_acks,
      return_reqs => accessMemory_return_reqs,
      return_acks => accessMemory_return_acks,
      call_data  => accessMemory_call_data,
      call_tag  => accessMemory_call_tag,
      return_tag  => accessMemory_return_tag,
      call_mtag => accessMemory_tag_in,
      return_mtag => accessMemory_tag_out,
      return_data =>accessMemory_return_data,
      call_mreq => accessMemory_start_req,
      call_mack => accessMemory_start_ack,
      return_mreq => accessMemory_fin_req,
      return_mack => accessMemory_fin_ack,
      call_mdata => accessMemory_in_args,
      return_mdata => accessMemory_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemory_instance:accessMemory-- 
    generic map(tag_length => 8)
    port map(-- 
      lock => accessMemory_lock,
      rwbar => accessMemory_rwbar,
      bmask => accessMemory_bmask,
      addr => accessMemory_addr,
      wdata => accessMemory_wdata,
      rdata => accessMemory_rdata,
      start_req => accessMemory_start_req,
      start_ack => accessMemory_start_ack,
      fin_req => accessMemory_fin_req,
      fin_ack => accessMemory_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemory_tag_in,
      tag_out => accessMemory_tag_out-- 
    ); -- 
  -- module acquireLock
  acquireLock_q_base_address <= acquireLock_in_args(35 downto 0);
  acquireLock_out_args <= acquireLock_m_ok ;
  -- call arbiter for module acquireLock
  acquireLock_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireLock_call_reqs,
      call_acks => acquireLock_call_acks,
      return_reqs => acquireLock_return_reqs,
      return_acks => acquireLock_return_acks,
      call_data  => acquireLock_call_data,
      call_tag  => acquireLock_call_tag,
      return_tag  => acquireLock_return_tag,
      call_mtag => acquireLock_tag_in,
      return_mtag => acquireLock_tag_out,
      return_data =>acquireLock_return_data,
      call_mreq => acquireLock_start_req,
      call_mack => acquireLock_start_ack,
      return_mreq => acquireLock_fin_req,
      return_mack => acquireLock_fin_ack,
      call_mdata => acquireLock_in_args,
      return_mdata => acquireLock_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireLock_instance:acquireLock-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => acquireLock_q_base_address,
      m_ok => acquireLock_m_ok,
      start_req => acquireLock_start_req,
      start_ack => acquireLock_start_ack,
      fin_req => acquireLock_fin_req,
      fin_ack => acquireLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(14 downto 14),
      accessMemory_call_acks => accessMemory_call_acks(14 downto 14),
      accessMemory_call_data => accessMemory_call_data(1649 downto 1540),
      accessMemory_call_tag => accessMemory_call_tag(44 downto 42),
      accessMemory_return_reqs => accessMemory_return_reqs(14 downto 14),
      accessMemory_return_acks => accessMemory_return_acks(14 downto 14),
      accessMemory_return_data => accessMemory_return_data(959 downto 896),
      accessMemory_return_tag => accessMemory_return_tag(44 downto 42),
      tag_in => acquireLock_tag_in,
      tag_out => acquireLock_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_q_base_address <= getQueueElement_in_args(67 downto 32);
  getQueueElement_read_index <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 68,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => getQueueElement_q_base_address,
      read_index => getQueueElement_read_index,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(11 downto 11),
      accessMemory_call_acks => accessMemory_call_acks(11 downto 11),
      accessMemory_call_data => accessMemory_call_data(1319 downto 1210),
      accessMemory_call_tag => accessMemory_call_tag(35 downto 33),
      accessMemory_return_reqs => accessMemory_return_reqs(11 downto 11),
      accessMemory_return_acks => accessMemory_return_acks(11 downto 11),
      accessMemory_return_data => accessMemory_return_data(767 downto 704),
      accessMemory_return_tag => accessMemory_return_tag(35 downto 33),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueueLength
  getQueueLength_q_base_address <= getQueueLength_in_args(35 downto 0);
  getQueueLength_out_args <= getQueueLength_Queue_Length ;
  -- call arbiter for module getQueueLength
  getQueueLength_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueLength_call_reqs,
      call_acks => getQueueLength_call_acks,
      return_reqs => getQueueLength_return_reqs,
      return_acks => getQueueLength_return_acks,
      call_data  => getQueueLength_call_data,
      call_tag  => getQueueLength_call_tag,
      return_tag  => getQueueLength_return_tag,
      call_mtag => getQueueLength_tag_in,
      return_mtag => getQueueLength_tag_out,
      return_data =>getQueueLength_return_data,
      call_mreq => getQueueLength_start_req,
      call_mack => getQueueLength_start_ack,
      return_mreq => getQueueLength_fin_req,
      return_mack => getQueueLength_fin_ack,
      call_mdata => getQueueLength_in_args,
      return_mdata => getQueueLength_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueLength_instance:getQueueLength-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueueLength_q_base_address,
      Queue_Length => getQueueLength_Queue_Length,
      start_req => getQueueLength_start_req,
      start_ack => getQueueLength_start_ack,
      fin_req => getQueueLength_fin_req,
      fin_ack => getQueueLength_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(7 downto 7),
      accessMemory_call_acks => accessMemory_call_acks(7 downto 7),
      accessMemory_call_data => accessMemory_call_data(879 downto 770),
      accessMemory_call_tag => accessMemory_call_tag(23 downto 21),
      accessMemory_return_reqs => accessMemory_return_reqs(7 downto 7),
      accessMemory_return_acks => accessMemory_return_acks(7 downto 7),
      accessMemory_return_data => accessMemory_return_data(511 downto 448),
      accessMemory_return_tag => accessMemory_return_tag(23 downto 21),
      tag_in => getQueueLength_tag_in,
      tag_out => getQueueLength_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_q_base_address <= getQueuePointers_in_args(35 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(8 downto 8),
      accessMemory_call_acks => accessMemory_call_acks(8 downto 8),
      accessMemory_call_data => accessMemory_call_data(989 downto 880),
      accessMemory_call_tag => accessMemory_call_tag(26 downto 24),
      accessMemory_return_reqs => accessMemory_return_reqs(8 downto 8),
      accessMemory_return_acks => accessMemory_return_acks(8 downto 8),
      accessMemory_return_data => accessMemory_return_data(575 downto 512),
      accessMemory_return_tag => accessMemory_return_tag(26 downto 24),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTotalMessages
  getTotalMessages_q_base_address <= getTotalMessages_in_args(35 downto 0);
  getTotalMessages_out_args <= getTotalMessages_total_msgs ;
  -- call arbiter for module getTotalMessages
  getTotalMessages_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTotalMessages_call_reqs,
      call_acks => getTotalMessages_call_acks,
      return_reqs => getTotalMessages_return_reqs,
      return_acks => getTotalMessages_return_acks,
      call_data  => getTotalMessages_call_data,
      call_tag  => getTotalMessages_call_tag,
      return_tag  => getTotalMessages_return_tag,
      call_mtag => getTotalMessages_tag_in,
      return_mtag => getTotalMessages_tag_out,
      return_data =>getTotalMessages_return_data,
      call_mreq => getTotalMessages_start_req,
      call_mack => getTotalMessages_start_ack,
      return_mreq => getTotalMessages_fin_req,
      return_mack => getTotalMessages_fin_ack,
      call_mdata => getTotalMessages_in_args,
      return_mdata => getTotalMessages_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTotalMessages_instance:getTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getTotalMessages_q_base_address,
      total_msgs => getTotalMessages_total_msgs,
      start_req => getTotalMessages_start_req,
      start_ack => getTotalMessages_start_ack,
      fin_req => getTotalMessages_fin_req,
      fin_ack => getTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(13 downto 13),
      accessMemory_call_acks => accessMemory_call_acks(13 downto 13),
      accessMemory_call_data => accessMemory_call_data(1539 downto 1430),
      accessMemory_call_tag => accessMemory_call_tag(41 downto 39),
      accessMemory_return_reqs => accessMemory_return_reqs(13 downto 13),
      accessMemory_return_acks => accessMemory_return_acks(13 downto 13),
      accessMemory_return_data => accessMemory_return_data(895 downto 832),
      accessMemory_return_tag => accessMemory_return_tag(41 downto 39),
      tag_in => getTotalMessages_tag_in,
      tag_out => getTotalMessages_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_queue_index <= getTxPacketPointerFromServer_in_args(5 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 33,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      queue_index => getTxPacketPointerFromServer_queue_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      AccessRegister_call_reqs => AccessRegister_call_reqs(2 downto 2),
      AccessRegister_call_acks => AccessRegister_call_acks(2 downto 2),
      AccessRegister_call_data => AccessRegister_call_data(128 downto 86),
      AccessRegister_call_tag => AccessRegister_call_tag(5 downto 4),
      AccessRegister_return_reqs => AccessRegister_return_reqs(2 downto 2),
      AccessRegister_return_acks => AccessRegister_return_acks(2 downto 2),
      AccessRegister_return_data => AccessRegister_return_data(95 downto 64),
      AccessRegister_return_tag => AccessRegister_return_tag(5 downto 4),
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(36 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(32 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(35 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(35 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(35 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(71 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(19 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(54 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(4 downto 3),
      AccessRegister_call_acks => AccessRegister_call_acks(4 downto 3),
      AccessRegister_call_data => AccessRegister_call_data(214 downto 129),
      AccessRegister_call_tag => AccessRegister_call_tag(9 downto 6),
      AccessRegister_return_reqs => AccessRegister_return_reqs(4 downto 3),
      AccessRegister_return_acks => AccessRegister_return_acks(4 downto 3),
      AccessRegister_return_data => AccessRegister_return_data(159 downto 96),
      AccessRegister_return_tag => AccessRegister_return_tag(9 downto 6),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module popFromQueue
  popFromQueue_lock <= popFromQueue_in_args(36 downto 36);
  popFromQueue_q_base_address <= popFromQueue_in_args(35 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 37,
      return_data_width => 33,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => popFromQueue_lock,
      q_base_address => popFromQueue_q_base_address,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(6 downto 6),
      accessMemory_call_acks => accessMemory_call_acks(6 downto 6),
      accessMemory_call_data => accessMemory_call_data(769 downto 660),
      accessMemory_call_tag => accessMemory_call_tag(20 downto 18),
      accessMemory_return_reqs => accessMemory_return_reqs(6 downto 6),
      accessMemory_return_acks => accessMemory_return_acks(6 downto 6),
      accessMemory_return_data => accessMemory_return_data(447 downto 384),
      accessMemory_return_tag => accessMemory_return_tag(20 downto 18),
      acquireLock_call_reqs => acquireLock_call_reqs(1 downto 1),
      acquireLock_call_acks => acquireLock_call_acks(1 downto 1),
      acquireLock_call_data => acquireLock_call_data(71 downto 36),
      acquireLock_call_tag => acquireLock_call_tag(1 downto 1),
      acquireLock_return_reqs => acquireLock_return_reqs(1 downto 1),
      acquireLock_return_acks => acquireLock_return_acks(1 downto 1),
      acquireLock_return_data => acquireLock_return_data(1 downto 1),
      acquireLock_return_tag => acquireLock_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 36),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      getQueueLength_call_reqs => getQueueLength_call_reqs(1 downto 1),
      getQueueLength_call_acks => getQueueLength_call_acks(1 downto 1),
      getQueueLength_call_data => getQueueLength_call_data(71 downto 36),
      getQueueLength_call_tag => getQueueLength_call_tag(1 downto 1),
      getQueueLength_return_reqs => getQueueLength_return_reqs(1 downto 1),
      getQueueLength_return_acks => getQueueLength_return_acks(1 downto 1),
      getQueueLength_return_data => getQueueLength_return_data(63 downto 32),
      getQueueLength_return_tag => getQueueLength_return_tag(1 downto 1),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(1 downto 1),
      getTotalMessages_call_acks => getTotalMessages_call_acks(1 downto 1),
      getTotalMessages_call_data => getTotalMessages_call_data(71 downto 36),
      getTotalMessages_call_tag => getTotalMessages_call_tag(1 downto 1),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(1 downto 1),
      getTotalMessages_return_acks => getTotalMessages_return_acks(1 downto 1),
      getTotalMessages_return_data => getTotalMessages_return_data(63 downto 32),
      getTotalMessages_return_tag => getTotalMessages_return_tag(1 downto 1),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(67 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(31 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(199 downto 100),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      updateTotalMessages_call_reqs => updateTotalMessages_call_reqs(1 downto 1),
      updateTotalMessages_call_acks => updateTotalMessages_call_acks(1 downto 1),
      updateTotalMessages_call_data => updateTotalMessages_call_data(135 downto 68),
      updateTotalMessages_call_tag => updateTotalMessages_call_tag(1 downto 1),
      updateTotalMessages_return_reqs => updateTotalMessages_return_reqs(1 downto 1),
      updateTotalMessages_return_acks => updateTotalMessages_return_acks(1 downto 1),
      updateTotalMessages_return_tag => updateTotalMessages_return_tag(1 downto 1),
      releaseLock_call_reqs => releaseLock_call_reqs(1 downto 1),
      releaseLock_call_acks => releaseLock_call_acks(1 downto 1),
      releaseLock_call_data => releaseLock_call_data(71 downto 36),
      releaseLock_call_tag => releaseLock_call_tag(1 downto 1),
      releaseLock_return_reqs => releaseLock_return_reqs(1 downto 1),
      releaseLock_return_acks => releaseLock_return_acks(1 downto 1),
      releaseLock_return_tag => releaseLock_return_tag(1 downto 1),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(35 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(11 downto 6),
      AccessRegister_call_reqs => AccessRegister_call_reqs(6 downto 6),
      AccessRegister_call_acks => AccessRegister_call_acks(6 downto 6),
      AccessRegister_call_data => AccessRegister_call_data(300 downto 258),
      AccessRegister_call_tag => AccessRegister_call_tag(13 downto 12),
      AccessRegister_return_reqs => AccessRegister_return_reqs(6 downto 6),
      AccessRegister_return_acks => AccessRegister_return_acks(6 downto 6),
      AccessRegister_return_data => AccessRegister_return_data(223 downto 192),
      AccessRegister_return_tag => AccessRegister_return_tag(13 downto 12),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(206 downto 138),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module pushIntoQueue
  pushIntoQueue_lock <= pushIntoQueue_in_args(68 downto 68);
  pushIntoQueue_q_base_address <= pushIntoQueue_in_args(67 downto 32);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(31 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 69,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => pushIntoQueue_lock,
      q_base_address => pushIntoQueue_q_base_address,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(4 downto 4),
      accessMemory_call_acks => accessMemory_call_acks(4 downto 4),
      accessMemory_call_data => accessMemory_call_data(549 downto 440),
      accessMemory_call_tag => accessMemory_call_tag(14 downto 12),
      accessMemory_return_reqs => accessMemory_return_reqs(4 downto 4),
      accessMemory_return_acks => accessMemory_return_acks(4 downto 4),
      accessMemory_return_data => accessMemory_return_data(319 downto 256),
      accessMemory_return_tag => accessMemory_return_tag(14 downto 12),
      acquireLock_call_reqs => acquireLock_call_reqs(0 downto 0),
      acquireLock_call_acks => acquireLock_call_acks(0 downto 0),
      acquireLock_call_data => acquireLock_call_data(35 downto 0),
      acquireLock_call_tag => acquireLock_call_tag(0 downto 0),
      acquireLock_return_reqs => acquireLock_return_reqs(0 downto 0),
      acquireLock_return_acks => acquireLock_return_acks(0 downto 0),
      acquireLock_return_data => acquireLock_return_data(0 downto 0),
      acquireLock_return_tag => acquireLock_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(35 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      getQueueLength_call_reqs => getQueueLength_call_reqs(0 downto 0),
      getQueueLength_call_acks => getQueueLength_call_acks(0 downto 0),
      getQueueLength_call_data => getQueueLength_call_data(35 downto 0),
      getQueueLength_call_tag => getQueueLength_call_tag(0 downto 0),
      getQueueLength_return_reqs => getQueueLength_return_reqs(0 downto 0),
      getQueueLength_return_acks => getQueueLength_return_acks(0 downto 0),
      getQueueLength_return_data => getQueueLength_return_data(31 downto 0),
      getQueueLength_return_tag => getQueueLength_return_tag(0 downto 0),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(0 downto 0),
      getTotalMessages_call_acks => getTotalMessages_call_acks(0 downto 0),
      getTotalMessages_call_data => getTotalMessages_call_data(35 downto 0),
      getTotalMessages_call_tag => getTotalMessages_call_tag(0 downto 0),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(0 downto 0),
      getTotalMessages_return_acks => getTotalMessages_return_acks(0 downto 0),
      getTotalMessages_return_data => getTotalMessages_return_data(31 downto 0),
      getTotalMessages_return_tag => getTotalMessages_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(99 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      updateTotalMessages_call_reqs => updateTotalMessages_call_reqs(0 downto 0),
      updateTotalMessages_call_acks => updateTotalMessages_call_acks(0 downto 0),
      updateTotalMessages_call_data => updateTotalMessages_call_data(67 downto 0),
      updateTotalMessages_call_tag => updateTotalMessages_call_tag(0 downto 0),
      updateTotalMessages_return_reqs => updateTotalMessages_return_reqs(0 downto 0),
      updateTotalMessages_return_acks => updateTotalMessages_return_acks(0 downto 0),
      updateTotalMessages_return_tag => updateTotalMessages_return_tag(0 downto 0),
      releaseLock_call_reqs => releaseLock_call_reqs(0 downto 0),
      releaseLock_call_acks => releaseLock_call_acks(0 downto 0),
      releaseLock_call_data => releaseLock_call_data(35 downto 0),
      releaseLock_call_tag => releaseLock_call_tag(0 downto 0),
      releaseLock_return_reqs => releaseLock_return_reqs(0 downto 0),
      releaseLock_return_acks => releaseLock_return_acks(0 downto 0),
      releaseLock_return_tag => releaseLock_return_tag(0 downto 0),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(99 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseLock
  releaseLock_q_base_address <= releaseLock_in_args(35 downto 0);
  -- call arbiter for module releaseLock
  releaseLock_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseLock_call_reqs,
      call_acks => releaseLock_call_acks,
      return_reqs => releaseLock_return_reqs,
      return_acks => releaseLock_return_acks,
      call_data  => releaseLock_call_data,
      call_tag  => releaseLock_call_tag,
      return_tag  => releaseLock_return_tag,
      call_mtag => releaseLock_tag_in,
      return_mtag => releaseLock_tag_out,
      call_mreq => releaseLock_start_req,
      call_mack => releaseLock_start_ack,
      return_mreq => releaseLock_fin_req,
      return_mack => releaseLock_fin_ack,
      call_mdata => releaseLock_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseLock_instance:releaseLock-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => releaseLock_q_base_address,
      start_req => releaseLock_start_req,
      start_ack => releaseLock_start_ack,
      fin_req => releaseLock_fin_req,
      fin_ack => releaseLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(10 downto 10),
      accessMemory_call_acks => accessMemory_call_acks(10 downto 10),
      accessMemory_call_data => accessMemory_call_data(1209 downto 1100),
      accessMemory_call_tag => accessMemory_call_tag(32 downto 30),
      accessMemory_return_reqs => accessMemory_return_reqs(10 downto 10),
      accessMemory_return_acks => accessMemory_return_acks(10 downto 10),
      accessMemory_return_data => accessMemory_return_data(703 downto 640),
      accessMemory_return_tag => accessMemory_return_tag(32 downto 30),
      tag_in => releaseLock_tag_in,
      tag_out => releaseLock_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_q_base_address <= setQueueElement_in_args(99 downto 64);
  setQueueElement_write_index <= setQueueElement_in_args(63 downto 32);
  setQueueElement_q_w_data <= setQueueElement_in_args(31 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 100,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => setQueueElement_q_base_address,
      write_index => setQueueElement_write_index,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(2 downto 2),
      accessMemory_call_acks => accessMemory_call_acks(2 downto 2),
      accessMemory_call_data => accessMemory_call_data(329 downto 220),
      accessMemory_call_tag => accessMemory_call_tag(8 downto 6),
      accessMemory_return_reqs => accessMemory_return_reqs(2 downto 2),
      accessMemory_return_acks => accessMemory_return_acks(2 downto 2),
      accessMemory_return_data => accessMemory_return_data(191 downto 128),
      accessMemory_return_tag => accessMemory_return_tag(8 downto 6),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_q_base_address <= setQueuePointers_in_args(99 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 100,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(15 downto 15),
      accessMemory_call_acks => accessMemory_call_acks(15 downto 15),
      accessMemory_call_data => accessMemory_call_data(1759 downto 1650),
      accessMemory_call_tag => accessMemory_call_tag(47 downto 45),
      accessMemory_return_reqs => accessMemory_return_reqs(15 downto 15),
      accessMemory_return_acks => accessMemory_return_acks(15 downto 15),
      accessMemory_return_data => accessMemory_return_data(1023 downto 960),
      accessMemory_return_tag => accessMemory_return_tag(47 downto 45),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      FREE_Q => FREE_Q,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      CONTROL_REGISTER => CONTROL_REGISTER,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(1 downto 1),
      AccessRegister_call_acks => AccessRegister_call_acks(1 downto 1),
      AccessRegister_call_data => AccessRegister_call_data(85 downto 43),
      AccessRegister_call_tag => AccessRegister_call_tag(3 downto 2),
      AccessRegister_return_reqs => AccessRegister_return_reqs(1 downto 1),
      AccessRegister_return_acks => AccessRegister_return_acks(1 downto 1),
      AccessRegister_return_data => AccessRegister_return_data(63 downto 32),
      AccessRegister_return_tag => AccessRegister_return_tag(3 downto 2),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(68 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(5 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(32 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(31 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_packet_pointer <= transmitPacket_in_args(31 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(0 downto 0),
      AccessRegister_call_acks => AccessRegister_call_acks(0 downto 0),
      AccessRegister_call_data => AccessRegister_call_data(42 downto 0),
      AccessRegister_call_tag => AccessRegister_call_tag(1 downto 0),
      AccessRegister_return_reqs => AccessRegister_return_reqs(0 downto 0),
      AccessRegister_return_acks => AccessRegister_return_acks(0 downto 0),
      AccessRegister_return_data => AccessRegister_return_data(31 downto 0),
      AccessRegister_return_tag => AccessRegister_return_tag(1 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(1 downto 0),
      accessMemory_call_acks => accessMemory_call_acks(1 downto 0),
      accessMemory_call_data => accessMemory_call_data(219 downto 0),
      accessMemory_call_tag => accessMemory_call_tag(5 downto 0),
      accessMemory_return_reqs => accessMemory_return_reqs(1 downto 0),
      accessMemory_return_acks => accessMemory_return_acks(1 downto 0),
      accessMemory_return_data => accessMemory_return_data(127 downto 0),
      accessMemory_return_tag => accessMemory_return_tag(5 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module updateTotalMessages
  updateTotalMessages_q_base_address <= updateTotalMessages_in_args(67 downto 32);
  updateTotalMessages_updated_total_msgs <= updateTotalMessages_in_args(31 downto 0);
  -- call arbiter for module updateTotalMessages
  updateTotalMessages_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 68,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => updateTotalMessages_call_reqs,
      call_acks => updateTotalMessages_call_acks,
      return_reqs => updateTotalMessages_return_reqs,
      return_acks => updateTotalMessages_return_acks,
      call_data  => updateTotalMessages_call_data,
      call_tag  => updateTotalMessages_call_tag,
      return_tag  => updateTotalMessages_return_tag,
      call_mtag => updateTotalMessages_tag_in,
      return_mtag => updateTotalMessages_tag_out,
      call_mreq => updateTotalMessages_start_req,
      call_mack => updateTotalMessages_start_ack,
      return_mreq => updateTotalMessages_fin_req,
      return_mack => updateTotalMessages_fin_ack,
      call_mdata => updateTotalMessages_in_args,
      clk => clk, 
      reset => reset --
    ); --
  updateTotalMessages_instance:updateTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => updateTotalMessages_q_base_address,
      updated_total_msgs => updateTotalMessages_updated_total_msgs,
      start_req => updateTotalMessages_start_req,
      start_ack => updateTotalMessages_start_ack,
      fin_req => updateTotalMessages_fin_req,
      fin_ack => updateTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(9 downto 9),
      accessMemory_call_acks => accessMemory_call_acks(9 downto 9),
      accessMemory_call_data => accessMemory_call_data(1099 downto 990),
      accessMemory_call_tag => accessMemory_call_tag(29 downto 27),
      accessMemory_return_reqs => accessMemory_return_reqs(9 downto 9),
      accessMemory_return_acks => accessMemory_return_acks(9 downto 9),
      accessMemory_return_data => accessMemory_return_data(639 downto 576),
      accessMemory_return_tag => accessMemory_return_tag(29 downto 27),
      tag_in => updateTotalMessages_tag_in,
      tag_out => updateTotalMessages_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(54 downto 19);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(18 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 55,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(3 downto 3),
      accessMemory_call_acks => accessMemory_call_acks(3 downto 3),
      accessMemory_call_data => accessMemory_call_data(439 downto 330),
      accessMemory_call_tag => accessMemory_call_tag(11 downto 9),
      accessMemory_return_reqs => accessMemory_return_reqs(3 downto 3),
      accessMemory_return_acks => accessMemory_return_acks(3 downto 3),
      accessMemory_return_data => accessMemory_return_data(255 downto 192),
      accessMemory_return_tag => accessMemory_return_tag(11 downto 9),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(35 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_buf_position_out ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      buf_position_out => writeEthernetHeaderToMem_buf_position_out,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(5 downto 5),
      accessMemory_call_acks => accessMemory_call_acks(5 downto 5),
      accessMemory_call_data => accessMemory_call_data(659 downto 550),
      accessMemory_call_tag => accessMemory_call_tag(17 downto 15),
      accessMemory_return_reqs => accessMemory_return_reqs(5 downto 5),
      accessMemory_return_acks => accessMemory_return_acks(5 downto 5),
      accessMemory_return_data => accessMemory_return_data(383 downto 320),
      accessMemory_return_tag => accessMemory_return_tag(17 downto 15),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(71 downto 36);
  writePayloadToMem_buf_pointer <= writePayloadToMem_in_args(35 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_32 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 20,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      buf_pointer => writePayloadToMem_buf_pointer,
      packet_size_32 => writePayloadToMem_packet_size_32,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(12 downto 12),
      accessMemory_call_acks => accessMemory_call_acks(12 downto 12),
      accessMemory_call_data => accessMemory_call_data(1429 downto 1320),
      accessMemory_call_tag => accessMemory_call_tag(38 downto 36),
      accessMemory_return_reqs => accessMemory_return_reqs(12 downto 12),
      accessMemory_return_acks => accessMemory_return_acks(12 downto 12),
      accessMemory_return_data => accessMemory_return_data(831 downto 768),
      accessMemory_return_tag => accessMemory_return_tag(38 downto 36),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => CONTROL_REGISTER,
      write_req => CONTROL_REGISTER_pipe_write_req,
      write_ack => CONTROL_REGISTER_pipe_write_ack,
      write_data => CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  FREE_Q_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe FREE_Q",
      volatile_flag => false,
      num_writes => 1,
      data_width => 36 --
    ) 
    port map( -- 
      read_data => FREE_Q,
      write_req => FREE_Q_pipe_write_req,
      write_ack => FREE_Q_pipe_write_ack,
      write_data => FREE_Q_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MAC_ENABLE_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe MAC_ENABLE",
      volatile_flag => false,
      num_writes => 1,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => MAC_ENABLE,
      write_req => MAC_ENABLE_pipe_write_req,
      write_ack => MAC_ENABLE_pipe_write_ack,
      write_data => MAC_ENABLE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_REQUEST_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_REQUEST_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 43,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_RESPONSE_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => NUMBER_OF_SERVERS,
      write_req => NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  enable_mac_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe enable_mac",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => enable_mac_pipe_read_req,
      read_ack => enable_mac_pipe_read_ack,
      read_data => enable_mac_pipe_read_data,
      write_req => enable_mac_pipe_write_req,
      write_ack => enable_mac_pipe_write_ack,
      write_data => enable_mac_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 2,
      addr_width => 6,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;


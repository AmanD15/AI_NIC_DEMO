-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_mac_bridge_lib;
use nic_mac_bridge_lib.rx_concat_system_global_package.all;
entity rx_concat is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_in_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    rx_in_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    rx_in_pipe_pipe_read_data : in   std_logic_vector(9 downto 0);
    rx_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    rx_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    rx_out_pipe_pipe_write_data : out  std_logic_vector(72 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity rx_concat;
architecture rx_concat_arch of rx_concat is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal rx_concat_CP_3_start: Boolean;
  signal rx_concat_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_9_branch_req_0 : boolean;
  signal phi_stmt_11_req_0 : boolean;
  signal phi_stmt_11_ack_0 : boolean;
  signal phi_stmt_11_req_1 : boolean;
  signal next_CIRCULANT_137_26_buf_req_0 : boolean;
  signal next_CIRCULANT_137_26_buf_ack_0 : boolean;
  signal next_CIRCULANT_137_26_buf_req_1 : boolean;
  signal next_CIRCULANT_137_26_buf_ack_1 : boolean;
  signal RPIPE_rx_in_pipe_29_inst_req_0 : boolean;
  signal RPIPE_rx_in_pipe_29_inst_ack_0 : boolean;
  signal RPIPE_rx_in_pipe_29_inst_req_1 : boolean;
  signal RPIPE_rx_in_pipe_29_inst_ack_1 : boolean;
  signal WPIPE_rx_out_pipe_146_inst_req_0 : boolean;
  signal WPIPE_rx_out_pipe_146_inst_ack_0 : boolean;
  signal WPIPE_rx_out_pipe_146_inst_req_1 : boolean;
  signal WPIPE_rx_out_pipe_146_inst_ack_1 : boolean;
  signal do_while_stmt_9_branch_ack_0 : boolean;
  signal do_while_stmt_9_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "rx_concat_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  rx_concat_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "rx_concat_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_concat_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= rx_concat_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_concat_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  rx_concat_CP_3: Block -- control-path 
    signal rx_concat_CP_3_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    rx_concat_CP_3_elements(0) <= rx_concat_CP_3_start;
    rx_concat_CP_3_symbol <= rx_concat_CP_3_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_8/$entry
      -- CP-element group 0: 	 branch_block_stmt_8/branch_block_stmt_8__entry__
      -- CP-element group 0: 	 branch_block_stmt_8/do_while_stmt_9__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	45 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_8/$exit
      -- CP-element group 1: 	 branch_block_stmt_8/branch_block_stmt_8__exit__
      -- CP-element group 1: 	 branch_block_stmt_8/do_while_stmt_9__exit__
      -- 
    rx_concat_CP_3_elements(1) <= rx_concat_CP_3_elements(45);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_8/do_while_stmt_9/$entry
      -- CP-element group 2: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9__entry__
      -- 
    rx_concat_CP_3_elements(2) <= rx_concat_CP_3_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	45 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9__exit__
      -- 
    -- Element group rx_concat_CP_3_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_8/do_while_stmt_9/loop_back
      -- 
    -- Element group rx_concat_CP_3_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	43 
    -- CP-element group 5: 	44 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_8/do_while_stmt_9/condition_done
      -- CP-element group 5: 	 branch_block_stmt_8/do_while_stmt_9/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_8/do_while_stmt_9/loop_taken/$entry
      -- 
    rx_concat_CP_3_elements(5) <= rx_concat_CP_3_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	42 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_8/do_while_stmt_9/loop_body_done
      -- 
    rx_concat_CP_3_elements(6) <= rx_concat_CP_3_elements(42);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/back_edge_to_loop_body
      -- 
    rx_concat_CP_3_elements(7) <= rx_concat_CP_3_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/first_time_through_loop_body
      -- 
    rx_concat_CP_3_elements(8) <= rx_concat_CP_3_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	41 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_27_sample_start_
      -- 
    -- Element group rx_concat_CP_3_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	41 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/condition_evaluated
      -- 
    condition_evaluated_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(10), ack => do_while_stmt_9_branch_req_0); -- 
    rx_concat_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(15) & rx_concat_CP_3_elements(41);
      gj_rx_concat_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	16 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_sample_start__ps
      -- 
    rx_concat_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(9) & rx_concat_CP_3_elements(16) & rx_concat_CP_3_elements(15);
      gj_rx_concat_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	36 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	42 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_27_sample_completed_
      -- 
    rx_concat_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(18) & rx_concat_CP_3_elements(36);
      gj_rx_concat_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	42 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group rx_concat_CP_3_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => rx_concat_CP_3_elements(12), ack => rx_concat_CP_3_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	33 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	35 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/aggregated_phi_update_req
      -- CP-element group 14: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_update_start__ps
      -- 
    rx_concat_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(17) & rx_concat_CP_3_elements(33);
      gj_rx_concat_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	37 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/aggregated_phi_update_ack
      -- 
    rx_concat_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(19) & rx_concat_CP_3_elements(37);
      gj_rx_concat_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_sample_start_
      -- 
    rx_concat_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(9) & rx_concat_CP_3_elements(12);
      gj_rx_concat_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	39 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_update_start_
      -- 
    rx_concat_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(9) & rx_concat_CP_3_elements(39);
      gj_rx_concat_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18: 	35 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_sample_completed__ps
      -- 
    -- Element group rx_concat_CP_3_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	38 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_update_completed__ps
      -- 
    -- Element group rx_concat_CP_3_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_loopback_trigger
      -- 
    rx_concat_CP_3_elements(20) <= rx_concat_CP_3_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_loopback_sample_req
      -- CP-element group 21: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_loopback_sample_req_ps
      -- 
    phi_stmt_11_loopback_sample_req_43_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_11_loopback_sample_req_43_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(21), ack => phi_stmt_11_req_1); -- 
    -- Element group rx_concat_CP_3_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_entry_trigger
      -- 
    rx_concat_CP_3_elements(22) <= rx_concat_CP_3_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_entry_sample_req
      -- CP-element group 23: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_entry_sample_req_ps
      -- 
    phi_stmt_11_entry_sample_req_46_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_11_entry_sample_req_46_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(23), ack => phi_stmt_11_req_0); -- 
    -- Element group rx_concat_CP_3_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_phi_mux_ack
      -- CP-element group 24: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_11_phi_mux_ack_ps
      -- 
    phi_stmt_11_phi_mux_ack_49_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_11_ack_0, ack => rx_concat_CP_3_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_sample_completed_
      -- 
    -- Element group rx_concat_CP_3_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_update_start_
      -- 
    -- Element group rx_concat_CP_3_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_update_completed__ps
      -- 
    rx_concat_CP_3_elements(27) <= rx_concat_CP_3_elements(28);
    -- CP-element group 28:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	27 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/CONCAT_u68_u76_24_update_completed_
      -- 
    -- Element group rx_concat_CP_3_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => rx_concat_CP_3_elements(26), ack => rx_concat_CP_3_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Sample/req
      -- 
    req_70_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_70_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(29), ack => next_CIRCULANT_137_26_buf_req_0); -- 
    -- Element group rx_concat_CP_3_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_update_start_
      -- CP-element group 30: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Update/req
      -- 
    req_75_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_75_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(30), ack => next_CIRCULANT_137_26_buf_req_1); -- 
    -- Element group rx_concat_CP_3_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Sample/ack
      -- 
    ack_71_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_CIRCULANT_137_26_buf_ack_0, ack => rx_concat_CP_3_elements(31)); -- 
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/R_next_CIRCULANT_26_Update/ack
      -- 
    ack_76_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_CIRCULANT_137_26_buf_ack_1, ack => rx_concat_CP_3_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	39 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	14 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_27_update_start_
      -- 
    rx_concat_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(9) & rx_concat_CP_3_elements(39);
      gj_rx_concat_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Sample/rr
      -- 
    rr_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(34), ack => RPIPE_rx_in_pipe_29_inst_req_0); -- 
    rx_concat_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(11) & rx_concat_CP_3_elements(37);
      gj_rx_concat_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	14 
    -- CP-element group 35: 	18 
    -- CP-element group 35: 	36 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_update_start_
      -- CP-element group 35: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Update/cr
      -- 
    cr_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(35), ack => RPIPE_rx_in_pipe_29_inst_req_1); -- 
    rx_concat_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(14) & rx_concat_CP_3_elements(18) & rx_concat_CP_3_elements(36);
      gj_rx_concat_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: 	35 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Sample/ra
      -- 
    ra_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_rx_in_pipe_29_inst_ack_0, ack => rx_concat_CP_3_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	15 
    -- CP-element group 37: 	38 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	34 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/phi_stmt_27_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/RPIPE_rx_in_pipe_29_Update/ca
      -- 
    ca_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_rx_in_pipe_29_inst_ack_1, ack => rx_concat_CP_3_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	19 
    -- CP-element group 38: 	37 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Sample/req
      -- 
    req_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(38), ack => WPIPE_rx_out_pipe_146_inst_req_0); -- 
    rx_concat_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(19) & rx_concat_CP_3_elements(37) & rx_concat_CP_3_elements(40);
      gj_rx_concat_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	17 
    -- CP-element group 39: 	33 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_update_start_
      -- CP-element group 39: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Update/req
      -- 
    ack_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_rx_out_pipe_146_inst_ack_0, ack => rx_concat_CP_3_elements(39)); -- 
    req_108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => rx_concat_CP_3_elements(39), ack => WPIPE_rx_out_pipe_146_inst_req_1); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/WPIPE_rx_out_pipe_146_Update/ack
      -- 
    ack_109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_rx_out_pipe_146_inst_ack_1, ack => rx_concat_CP_3_elements(40)); -- 
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	9 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	10 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group rx_concat_CP_3_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => rx_concat_CP_3_elements(9), ack => rx_concat_CP_3_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	12 
    -- CP-element group 42: 	13 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	6 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_8/do_while_stmt_9/do_while_stmt_9_loop_body/$exit
      -- 
    rx_concat_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "rx_concat_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= rx_concat_CP_3_elements(12) & rx_concat_CP_3_elements(13) & rx_concat_CP_3_elements(40);
      gj_rx_concat_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => rx_concat_CP_3_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_8/do_while_stmt_9/loop_exit/$exit
      -- CP-element group 43: 	 branch_block_stmt_8/do_while_stmt_9/loop_exit/ack
      -- 
    ack_114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_9_branch_ack_0, ack => rx_concat_CP_3_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	5 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_8/do_while_stmt_9/loop_taken/$exit
      -- CP-element group 44: 	 branch_block_stmt_8/do_while_stmt_9/loop_taken/ack
      -- 
    ack_118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_9_branch_ack_1, ack => rx_concat_CP_3_elements(44)); -- 
    -- CP-element group 45:  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	3 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	1 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_8/do_while_stmt_9/$exit
      -- 
    rx_concat_CP_3_elements(45) <= rx_concat_CP_3_elements(3);
    rx_concat_do_while_stmt_9_terminator_119: loop_terminator -- 
      generic map (name => " rx_concat_do_while_stmt_9_terminator_119", max_iterations_in_flight =>7) 
      port map(loop_body_exit => rx_concat_CP_3_elements(6),loop_continue => rx_concat_CP_3_elements(44),loop_terminate => rx_concat_CP_3_elements(43),loop_back => rx_concat_CP_3_elements(4),loop_exit => rx_concat_CP_3_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_11_phi_seq_77_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= rx_concat_CP_3_elements(22);
      rx_concat_CP_3_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= rx_concat_CP_3_elements(25);
      rx_concat_CP_3_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= rx_concat_CP_3_elements(27);
      rx_concat_CP_3_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= rx_concat_CP_3_elements(20);
      rx_concat_CP_3_elements(29)<= src_sample_reqs(1);
      src_sample_acks(1)  <= rx_concat_CP_3_elements(31);
      rx_concat_CP_3_elements(30)<= src_update_reqs(1);
      src_update_acks(1)  <= rx_concat_CP_3_elements(32);
      rx_concat_CP_3_elements(21) <= phi_mux_reqs(1);
      phi_stmt_11_phi_seq_77 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_11_phi_seq_77") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => rx_concat_CP_3_elements(11), 
          phi_sample_ack => rx_concat_CP_3_elements(18), 
          phi_update_req => rx_concat_CP_3_elements(14), 
          phi_update_ack => rx_concat_CP_3_elements(19), 
          phi_mux_ack => rx_concat_CP_3_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_28_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= rx_concat_CP_3_elements(7);
        preds(1)  <= rx_concat_CP_3_elements(8);
        entry_tmerge_28 : transition_merge -- 
          generic map(name => " entry_tmerge_28")
          port map (preds => preds, symbol_out => rx_concat_CP_3_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u4_u4_79_wire : std_logic_vector(3 downto 0);
    signal AND_u1_u1_108_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_119_wire : std_logic_vector(0 downto 0);
    signal CIRCULANT_11 : std_logic_vector(75 downto 0);
    signal CONCAT_u1_u65_141_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u4_u7_101_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u64_u68_134_wire : std_logic_vector(67 downto 0);
    signal CONCAT_u68_u76_24_wire_constant : std_logic_vector(75 downto 0);
    signal CONCAT_u7_u8_91_wire : std_logic_vector(7 downto 0);
    signal EQ_u4_u1_56_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_107_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_118_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_122_wire_constant : std_logic_vector(7 downto 0);
    signal RPIPE_rx_in_pipe_29_wire : std_logic_vector(9 downto 0);
    signal RX_27 : std_logic_vector(9 downto 0);
    signal SHL_u64_u64_112_wire : std_logic_vector(63 downto 0);
    signal SHL_u8_u8_128_wire : std_logic_vector(7 downto 0);
    signal SUB_u4_u4_126_wire : std_logic_vector(3 downto 0);
    signal SUB_u4_u4_97_wire : std_logic_vector(3 downto 0);
    signal byte_mask_to_pipe_130 : std_logic_vector(7 downto 0);
    signal collected_dword_34 : std_logic_vector(63 downto 0);
    signal data_to_pipe_114 : std_logic_vector(63 downto 0);
    signal dword_to_pipe_65 : std_logic_vector(63 downto 0);
    signal konst_124_wire_constant : std_logic_vector(3 downto 0);
    signal konst_150_wire_constant : std_logic_vector(0 downto 0);
    signal konst_55_wire_constant : std_logic_vector(3 downto 0);
    signal konst_78_wire_constant : std_logic_vector(3 downto 0);
    signal konst_95_wire_constant : std_logic_vector(3 downto 0);
    signal left_shift_amount_103 : std_logic_vector(63 downto 0);
    signal next_CIRCULANT_137 : std_logic_vector(75 downto 0);
    signal next_CIRCULANT_137_26_buffered : std_logic_vector(75 downto 0);
    signal next_collected_dword_72 : std_logic_vector(63 downto 0);
    signal next_running_byte_count_81 : std_logic_vector(3 downto 0);
    signal next_running_byte_mask_93 : std_logic_vector(7 downto 0);
    signal running_byte_count_38 : std_logic_vector(3 downto 0);
    signal running_byte_mask_42 : std_logic_vector(7 downto 0);
    signal rx_data_51 : std_logic_vector(7 downto 0);
    signal rx_last_47 : std_logic_vector(0 downto 0);
    signal send_to_pipe_58 : std_logic_vector(0 downto 0);
    signal slice_62_wire : std_logic_vector(55 downto 0);
    signal slice_88_wire : std_logic_vector(6 downto 0);
    signal to_pipe_144 : std_logic_vector(72 downto 0);
    signal type_cast_100_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_127_wire : std_logic_vector(7 downto 0);
    signal type_cast_69_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_76_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    CONCAT_u68_u76_24_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000100000001";
    NOT_u8_u8_122_wire_constant <= "11111111";
    konst_124_wire_constant <= "1000";
    konst_150_wire_constant <= "1";
    konst_55_wire_constant <= "1000";
    konst_78_wire_constant <= "0001";
    konst_95_wire_constant <= "1000";
    type_cast_100_wire_constant <= "000";
    type_cast_69_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_76_wire_constant <= "0001";
    type_cast_85_wire_constant <= "00000001";
    type_cast_90_wire_constant <= "1";
    phi_stmt_11: Block -- phi operator 
      signal idata: std_logic_vector(151 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= CONCAT_u68_u76_24_wire_constant & next_CIRCULANT_137_26_buffered;
      req <= phi_stmt_11_req_0 & phi_stmt_11_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_11",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 76) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_11_ack_0,
          idata => idata,
          odata => CIRCULANT_11,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_11
    -- flow-through select operator MUX_113_inst
    data_to_pipe_114 <= dword_to_pipe_65 when (AND_u1_u1_108_wire(0) /=  '0') else SHL_u64_u64_112_wire;
    -- flow-through select operator MUX_129_inst
    byte_mask_to_pipe_130 <= NOT_u8_u8_122_wire_constant when (AND_u1_u1_119_wire(0) /=  '0') else SHL_u8_u8_128_wire;
    -- flow-through select operator MUX_71_inst
    next_collected_dword_72 <= type_cast_69_wire_constant when (send_to_pipe_58(0) /=  '0') else dword_to_pipe_65;
    -- flow-through select operator MUX_80_inst
    next_running_byte_count_81 <= type_cast_76_wire_constant when (send_to_pipe_58(0) /=  '0') else ADD_u4_u4_79_wire;
    -- flow-through select operator MUX_92_inst
    next_running_byte_mask_93 <= type_cast_85_wire_constant when (send_to_pipe_58(0) /=  '0') else CONCAT_u7_u8_91_wire;
    -- flow-through slice operator slice_33_inst
    collected_dword_34 <= CIRCULANT_11(75 downto 12);
    -- flow-through slice operator slice_37_inst
    running_byte_count_38 <= CIRCULANT_11(11 downto 8);
    -- flow-through slice operator slice_41_inst
    running_byte_mask_42 <= CIRCULANT_11(7 downto 0);
    -- flow-through slice operator slice_46_inst
    rx_last_47 <= RX_27(9 downto 9);
    -- flow-through slice operator slice_50_inst
    rx_data_51 <= RX_27(8 downto 1);
    -- flow-through slice operator slice_62_inst
    slice_62_wire <= collected_dword_34(55 downto 0);
    -- flow-through slice operator slice_88_inst
    slice_88_wire <= running_byte_mask_42(6 downto 0);
    next_CIRCULANT_137_26_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_CIRCULANT_137_26_buf_req_0;
      next_CIRCULANT_137_26_buf_ack_0<= wack(0);
      rreq(0) <= next_CIRCULANT_137_26_buf_req_1;
      next_CIRCULANT_137_26_buf_ack_1<= rack(0);
      next_CIRCULANT_137_26_buf : InterlockBuffer generic map ( -- 
        name => "next_CIRCULANT_137_26_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 76,
        out_data_width => 76,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_CIRCULANT_137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_CIRCULANT_137_26_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_27
    process(RPIPE_rx_in_pipe_29_wire) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 9 downto 0) := RPIPE_rx_in_pipe_29_wire(9 downto 0);
      RX_27 <= tmp_var; -- 
    end process;
    -- interlock type_cast_102_inst
    process(CONCAT_u4_u7_101_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 6 downto 0) := CONCAT_u4_u7_101_wire(6 downto 0);
      left_shift_amount_103 <= tmp_var; -- 
    end process;
    -- interlock type_cast_127_inst
    process(SUB_u4_u4_126_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 3 downto 0) := SUB_u4_u4_126_wire(3 downto 0);
      type_cast_127_wire <= tmp_var; -- 
    end process;
    do_while_stmt_9_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_150_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_9_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_9_branch_req_0,
          ack0 => do_while_stmt_9_branch_ack_0,
          ack1 => do_while_stmt_9_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u4_u4_79_inst
    ADD_u4_u4_79_wire <= std_logic_vector(unsigned(running_byte_count_38) + unsigned(konst_78_wire_constant));
    -- flow through binary operator AND_u1_u1_108_inst
    AND_u1_u1_108_wire <= (send_to_pipe_58 and NOT_u1_u1_107_wire);
    -- flow through binary operator AND_u1_u1_119_inst
    AND_u1_u1_119_wire <= (send_to_pipe_58 and NOT_u1_u1_118_wire);
    -- flow through binary operator CONCAT_u1_u65_141_inst
    process(rx_last_47, data_to_pipe_114) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_last_47, data_to_pipe_114, tmp_var);
      CONCAT_u1_u65_141_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u4_u7_101_inst
    process(SUB_u4_u4_97_wire) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(SUB_u4_u4_97_wire, type_cast_100_wire_constant, tmp_var);
      CONCAT_u4_u7_101_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u56_u64_64_inst
    process(slice_62_wire, rx_data_51) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_62_wire, rx_data_51, tmp_var);
      dword_to_pipe_65 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u64_u68_134_inst
    process(next_collected_dword_72, next_running_byte_count_81) -- 
      variable tmp_var : std_logic_vector(67 downto 0); -- 
    begin -- 
      ApConcat_proc(next_collected_dword_72, next_running_byte_count_81, tmp_var);
      CONCAT_u64_u68_134_wire <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u65_u73_143_inst
    process(CONCAT_u1_u65_141_wire, byte_mask_to_pipe_130) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u65_141_wire, byte_mask_to_pipe_130, tmp_var);
      to_pipe_144 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u68_u76_136_inst
    process(CONCAT_u64_u68_134_wire, next_running_byte_mask_93) -- 
      variable tmp_var : std_logic_vector(75 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u64_u68_134_wire, next_running_byte_mask_93, tmp_var);
      next_CIRCULANT_137 <= tmp_var; --
    end process;
    -- flow through binary operator CONCAT_u7_u8_91_inst
    process(slice_88_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_88_wire, type_cast_90_wire_constant, tmp_var);
      CONCAT_u7_u8_91_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u4_u1_56_inst
    process(running_byte_count_38) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(running_byte_count_38, konst_55_wire_constant, tmp_var);
      EQ_u4_u1_56_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_107_inst
    process(rx_last_47) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rx_last_47, tmp_var);
      NOT_u1_u1_107_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_118_inst
    process(rx_last_47) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rx_last_47, tmp_var);
      NOT_u1_u1_118_wire <= tmp_var; -- 
    end process;
    -- flow through binary operator OR_u1_u1_57_inst
    send_to_pipe_58 <= (rx_last_47 or EQ_u4_u1_56_wire);
    -- flow through binary operator SHL_u64_u64_112_inst
    process(dword_to_pipe_65, left_shift_amount_103) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(dword_to_pipe_65, left_shift_amount_103, tmp_var);
      SHL_u64_u64_112_wire <= tmp_var; --
    end process;
    -- flow through binary operator SHL_u8_u8_128_inst
    process(running_byte_mask_42, type_cast_127_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(running_byte_mask_42, type_cast_127_wire, tmp_var);
      SHL_u8_u8_128_wire <= tmp_var; --
    end process;
    -- flow through binary operator SUB_u4_u4_126_inst
    SUB_u4_u4_126_wire <= std_logic_vector(unsigned(konst_124_wire_constant) - unsigned(running_byte_count_38));
    -- flow through binary operator SUB_u4_u4_97_inst
    SUB_u4_u4_97_wire <= std_logic_vector(unsigned(konst_95_wire_constant) - unsigned(running_byte_count_38));
    -- shared inport operator group (0) : RPIPE_rx_in_pipe_29_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(9 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_rx_in_pipe_29_inst_req_0;
      RPIPE_rx_in_pipe_29_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_rx_in_pipe_29_inst_req_1;
      RPIPE_rx_in_pipe_29_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_rx_in_pipe_29_wire <= data_out(9 downto 0);
      rx_in_pipe_read_0_gI: SplitGuardInterface generic map(name => "rx_in_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      rx_in_pipe_read_0: InputPortRevised -- 
        generic map ( name => "rx_in_pipe_read_0", data_width => 10,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => rx_in_pipe_pipe_read_req(0),
          oack => rx_in_pipe_pipe_read_ack(0),
          odata => rx_in_pipe_pipe_read_data(9 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_rx_out_pipe_146_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_rx_out_pipe_146_inst_req_0;
      WPIPE_rx_out_pipe_146_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_rx_out_pipe_146_inst_req_1;
      WPIPE_rx_out_pipe_146_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_pipe_58(0);
      data_in <= to_pipe_144;
      rx_out_pipe_write_0_gI: SplitGuardInterface generic map(name => "rx_out_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      rx_out_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "rx_out_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => rx_out_pipe_pipe_write_req(0),
          oack => rx_out_pipe_pipe_write_ack(0),
          odata => rx_out_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end rx_concat_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library nic_mac_bridge_lib;
use nic_mac_bridge_lib.rx_concat_system_global_package.all;
entity rx_concat_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    rx_in_pipe_pipe_write_data: in std_logic_vector(9 downto 0);
    rx_in_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    rx_in_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    rx_out_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    rx_out_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    rx_out_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture rx_concat_system_arch  of rx_concat_system is -- system-architecture 
  -- declarations related to module rx_concat
  component rx_concat is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_in_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      rx_in_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rx_in_pipe_pipe_read_data : in   std_logic_vector(9 downto 0);
      rx_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      rx_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      rx_out_pipe_pipe_write_data : out  std_logic_vector(72 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module rx_concat
  signal rx_concat_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal rx_concat_tag_out   : std_logic_vector(1 downto 0);
  signal rx_concat_start_req : std_logic;
  signal rx_concat_start_ack : std_logic;
  signal rx_concat_fin_req   : std_logic;
  signal rx_concat_fin_ack : std_logic;
  -- aggregate signals for read from pipe rx_in_pipe
  signal rx_in_pipe_pipe_read_data: std_logic_vector(9 downto 0);
  signal rx_in_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal rx_in_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe rx_out_pipe
  signal rx_out_pipe_pipe_write_data: std_logic_vector(72 downto 0);
  signal rx_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal rx_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module rx_concat
  rx_concat_instance:rx_concat-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => rx_concat_start_req,
      start_ack => rx_concat_start_ack,
      fin_req => rx_concat_fin_req,
      fin_ack => rx_concat_fin_ack,
      clk => clk,
      reset => reset,
      rx_in_pipe_pipe_read_req => rx_in_pipe_pipe_read_req(0 downto 0),
      rx_in_pipe_pipe_read_ack => rx_in_pipe_pipe_read_ack(0 downto 0),
      rx_in_pipe_pipe_read_data => rx_in_pipe_pipe_read_data(9 downto 0),
      rx_out_pipe_pipe_write_req => rx_out_pipe_pipe_write_req(0 downto 0),
      rx_out_pipe_pipe_write_ack => rx_out_pipe_pipe_write_ack(0 downto 0),
      rx_out_pipe_pipe_write_data => rx_out_pipe_pipe_write_data(72 downto 0),
      tag_in => rx_concat_tag_in,
      tag_out => rx_concat_tag_out-- 
    ); -- 
  -- module will be run forever 
  rx_concat_tag_in <= (others => '0');
  rx_concat_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => rx_concat_start_req, start_ack => rx_concat_start_ack,  fin_req => rx_concat_fin_req,  fin_ack => rx_concat_fin_ack);
  rx_in_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe rx_in_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 10,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => rx_in_pipe_pipe_read_req,
      read_ack => rx_in_pipe_pipe_read_ack,
      read_data => rx_in_pipe_pipe_read_data,
      write_req => rx_in_pipe_pipe_write_req,
      write_ack => rx_in_pipe_pipe_write_ack,
      write_data => rx_in_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  rx_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe rx_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => rx_out_pipe_pipe_read_req,
      read_ack => rx_out_pipe_pipe_read_ack,
      read_data => rx_out_pipe_pipe_read_data,
      write_req => rx_out_pipe_pipe_write_req,
      write_ack => rx_out_pipe_pipe_write_ack,
      write_data => rx_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  -- 
end rx_concat_system_arch;



`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N0hMcXbI5hCFMXvbzZaWNMXky7Cb78UlPrOh26mC4IyomLPXkDt4pohvBi74RwhMjj/Bp6A1/EjU
BW4AL9d6yw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O4cgU289ETKimPPpC1lQoWfngvpNmR5tUZAEw+00K8UK2gEeqXn1hb3g7AZENGEwMii7hns4XQy8
DXQ5xw0Yp1Lt5kPvabj5mKM1bMdX8dvR9NHP3g1Qjd7okAVBl07/JG0NTnpHDOfWPgdIKiG5gomz
/inOtmJ9dyw3SQwornQ=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DU+IJVy0UCp9Ru4O1AHH4hAsURQvG4KWjfdJuBdXBn/Aw7vf76lLrDggWEsh/tDsD2w8gcTI1KZj
gte8Qz0RBjJA/tV/Q7C3IGP9sKs04WbpHeToWiLkJhGVSOi1cfBwcXqun7kk3rw8tbtRvnn4LLnQ
VVSnOUM0P3u3t9b+354=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VU2OWBPAFdMWY9YsdLW9vHBQultKfSyqJgSm8GFxf210g4AV7503RY1sTzcwbpKduWx2mEapVrlR
2+Drhdzv1Rts/cH1vI36ZrlUVzIXAPfly2Vw/ZI3vZ8ecksIx4K68q0S13FJLdHLryPXLuFGokYw
gCOZnAxTuOQQMCgsJA0iDJVXFdmLXzqwRYBXguqf1r+OMVPXs57gcwlgVB8r2wrtRxBvH0uRcmEd
9XDbIcnUXETCLhyRgVVpblWBh8bZbcQBY/zZZ/sbyAPD6J7Rp8CEPhLVVCsK4EjNey5PsDgo/izg
h4bUKLC5eF2W7tVckgp7jyOfw3DgIr/wn7RxeQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V2G0fgDEE2OFe05Cx8OR1KsgdINzVEXBIBadpSnPXIoTc7xRwAe4/VP6V+6MXz0QrLZuQHVAj7G3
9F/ijf7v4vM07B7zCCzqKWXPOd8bPZE51/A2H7Mt+ilGqjbh/VKLmxGs4hilsENWISKVXeBdKnPY
gj2HGvaphMJpBpJwjPAKBmbUyTX5Sd9nNIMzcSRJNulwiaiEOrABFlrZOI+c7bZY5sHmVeOtg9CQ
vhwpJiZDt2xEUYZdJ+nAzC0+NS9jg6KFWoyyUeNOwHZC9//fhh1MCUzJ0nZg2R4hBpRaxLZstp3w
PM0at5MBtCkDuhRItVUmq9A0HtCUCEmB412P1w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RN/6I+vbSUSbgQKZutSOM516q9s9JryaK6V/qqxo3gcYd+gU9W/srRAx8TWXTu0WbgzNnJ4y7Myb
hqdFZXcfJ/PxMgXPrrBTM9dc9q6Om0xxWrgSNxYalV3KY2vgAYOZai6mnccqhDfT+ZicibnnsYmh
yf5l9IBMwTbxQ9cpGytJTrr0jtjFG8izeH9CEj3vxYZQ4tA0TFJhsFvQhk2xXEnWnEBhTQbSX/B3
CADhGzXitOUqpBt3ylEkYkNM5wRAzze9LtBQhOCFWc4AJq4+3/P22qqco2g+VSDFNt7Sbc/BGwyj
q/3tdC0FZkEZB5DXnSDvgc9OVq2Fggic0aDyNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
iaxYaaoY/5xTFt2c8M0tGlrXM4N/DM5yeuEibfkumBAtVIC7iAa7xWJt8/5rQDlwIN5ywa11wy6G
GhBjDNeTFaFKIB2rr7Fl4tMwltZXdqJqhI0tN4Edm7gKZndbjiAQYtW21kCUeFhAZ+AlQnCDDpT+
jxcmgVQS2sLbZ3F0ud8OJNKpGktcgoXZWNss3tlknLzZro6/DZj9RrPutnuw5sEfz6xxFVdozrc5
tusWh76JQgz6u7g/pFOebhHGMNIHXun6iaIkaZGqx/LdNWvzg4RbNuwPFg21+jeh9vi1CRnzBuvf
f+/nz+S3sMnZND4fpp5g44AAjJF+PoWAZ49cqLEDsq9exu9q8JtQGsNdbR2z3T6pOmXvkyHaVh+r
aRm6UiyldFs4WDXtHLtEY62K8GgsLyYWlRxtrgJDHpCKCL5ub8ojJF2kTRT2aarND4e5PflYZYjp
3ym5ReincLUsmlhaf1+p730yJUMPMxK7u7KsOQ47f8f2iX62jshiYbm869wWLhjLzqGj0TD5QP1p
ptuLkp5C3Iqx3qNTRKG6FNtWlWjzg8zEBpfVhenjZopd1hZ9A5Ve0e6RkE5/s6tqvYNGbhLO+WHD
JfOvUncsiCZtcFlYhkKazEFuU7qe9zyyI+IILrppv2mrLU+R7fsUzUNIUy/GjaeowbSH/fGlHOUW
gRnbTwwdRzzMpFZQaV4z7LmQffvirV8bZ/2qXOgHIWLs/zRJZI9JBqens1jJliH9glQzuJ2MWaOf
wqwgFs0XDwoMJOhYqzm1ulDZ2rnpD1BwB2HBLkkdS2MQ0d2/g9Q/tt1A6wjE8uvXspevmEvCJUEa
XR8xSBKkVnj/mgZFYd2MWQsjX4q6X/pjDfXuXU2ucwC05e95Osm2AQ+7GVtsJL+0j70Znt80gAtn
bwhlPdWccyath2jJS/xMJsqzMKxE+y5nqtpzujRtKBIZTfJn4DJ3SMGlmp/khQaa/i9Jh0ei8pe6
HPhPor4KZ7wpYcGIOkBkRTelrI6WkL+IWXD4qsnDhm7UX3abV+JcnbympPUZ00BWFbRwBKf1t2OK
a0yd05QsUrUDs4VaD6Amb+f023x16VG5pEDWjW2QAbX5mzUsnDdcVWfkbd4uqgqKA4Q4F/6gSX0Z
zqw89bGR93RMrO6FVgpW3/U4pu92/BdccHzoG21PcW/uZJzcJPJsrL8HDCgTFhryKs/uWPU2wZig
ciScXrCC+7NNfpuz7ZIca2jKiDGD9Xs3nzmecSDRYJ0DqiRvELS+y+vfIxZQVD+zd/b3X1y6riGE
PjlI+2u5mMkYy2aZqoVtnF11wH7oxWKh4Hlr4ztx0Wu2vX7ShT13BP5KWLZ8FKd+jHIQEU6UQWIx
dq/ggHJck14ZTrXPSTSv3anZ7AZXMMdfGr1Sw7RcP1fbMndOY4lZGA8GBlcTPhh0PdpBW4Xn4dyU
mp6PN505BZWEBI1fZxwTnmwv9frbF/BZGvoFZBZVHPf32xwXrARku6Y4T+qe/o6juD84BiI8Bggz
d1hoMWj3i6lsHRh+UCtGIIX3C7/bCYzXdbcOoZcMe0m9iNx+vxY0m2/vSc6P15SOoeePoKMD0Fdf
M3JJoEZaImHs/mywXiT4hIOnNqeNKbMRIhR+gGvXNddi7ZtxLa4hyaWy7wRD5rt0B2CnEKksP4zT
OY2bcidFkA4JS05sA/38mXA1Z32I7I4skBPPuSZPOqn/9g/uMNqq5wm1rzGS2l0I4FVEaJ9631By
wqwhZB1t4P/7X8RhqYp9BT8WgNusJ83eTVeFEeHQs7ydd1F6XUCJsFwAVfRdIrJDBm/5FOvT6UxP
ZRGRa395tIlSiXVSvXkQOdPyij3rZa2qI06nptMMy8mtjXK4bxNxsoIF5LN03UKv+SSO9hMosPnt
DQ222sZSJCzcDA8Q7kpo0OBLHqjNaRK8BaYlW0473hnUIOCOxBASst8y8lfCdZZ84IepAQy5O44k
jzlcDS5mhXrhh88DUVp0g7YS0iSKC9CecC+5rf6iWvwrB7GdxzoG0w9y7QW22uYMYhUIjN+auubK
08hYL/lwbl9cMVjIpyx4pTQL/WP9+wG0Gp5GSHYLM9Cd1axesycaU4FkHTEmw68yZ1z5wUAhmvpZ
csHEIYxm31WKNvQYQe0WxnyUn3apBZkTMO8Pl9Dv8nYLYXQxrMdM0e/VjtQ1a58LO73sGmDrYXtm
+HIWdxKMgk3hV0NYwKV3vADJjwbfaCfzVREjnZNwpIAqIe+nHwD8Ywsxck4qzMTKZr7GVFIZfZiM
f+1h2OTs+CgAFi6NBE8jfWRaJem/wUknrD8BbhSkNNaTIDg+WPDboBgKKN1JggYDp+2b5ouJ1yU8
Aej1vAo0XG8B31ZQXEWidz74qWpCDQq25BPLb1ygTT70Bq6M0FNphffghQqoZZMImRu7XDa/2Y9d
5NxkibUW3yA2Uf7lNPkVyOv+mp74uI1/mcyTjAkEYAN7mKp+mZIf0rYof7ziNiUNvgxU1heegwla
vjOdv2LWCUbjeSHcpF2Yvhyg8AiUXEfTOYCBNmb1D0ffw6d1b66S0YQCu8cBwBtRJXClkjHrPkxJ
LHC614v6joK+F+CaX5EaMaqEolzfelgs94aLEh6bgiV5+jbzuS2EDn8UqEA3oFGhI9pOAh1JSWvX
IEkraMIAw8YPfy4Zi4gRp9sIs1HK2Hql2Dr163bh0d+N0EkEo/v1fD0DKXB+kC61Ov04YEjaoS0T
IS5CsuNRr5rG31JsJpQp2GeW4G1/I3AD/mVlje8ew5Rw7JDVxpRfT11fuvx5y3vd0AO8/OORNUYu
QFKAaWrIGdgf/PRPG/vMpCvl2OgCiNCdepEUolFIyQckLmh3luOyT12HJE1vUk9NfAcUpdqec66s
gTOi10CBdrmFNnAlWe1UUNJ81J9zSrJNM7rSANViDmXV2X6U/MydOCPzGf4AsKM2YknqPXSF3LGr
bFxlvpVzBvbx0Qb9aI4offggojkpQOL/Y2Bny8ZQnjGppk4wty48aATw/2rs3WqBkQQfRBQ7nnTl
m99h4T02yoIHg65TU8/qAkHQgf2NbxzdNtwzeTAH6odTuPO1+yZzLiK4nq39wn++U3mWqOQCQ9p/
UWr1VbWfL+WgAwIj70B2T8iCPbD3nLgfX4bHBD5ERDFMSa6S6pNoULekB14h/Y7c1n2M5F+iNFPz
VJ4xf404EqZBtQA3y5McYrjoIFxzvVmrxDkPMNt3FG7PpbJjCasyQ5mjPIsAcPfY576Qx2COhDAn
y76RqfTW34+BBUXeIFlSyowafuhg1ottRzUOlo4wc/8vVlLNDE+upAGes2T4i+LYMHjHu3UyzsAQ
mkgbJ7g/Y8x+u+pmP/8uxT1iAXjhRcQ5vP4FX4D39WFfvEn3sPKdDj+0YZoJ7oYljc0hapl8Tbo8
2XXsNdpKRA2wRWH4KnK1XqzXGrkex20wfdKPQDC75FDhtqcD4h2nkXgD9KCtneRuwK96+8Vveu6+
t8hgHveXW9pZAKTMOdEBpla/SmL+kpZIzOob1noxQgEmbRvlrGmcjubfDxHwdlxRu+PdwJJonZEN
LAoG1iymvuJhDwQEr0MQWZtXanhZhcCREvL9PHRtKgTRoQWNX4BtDZi9zXBBd+1fDnrjPZlwHVSy
aP/ke16Fn+969CpJr5foaw+xJupmyGa5qhTFmOkchi5BsQBCyIR4/z4SPB/EvCO6keGZmgdcYsOx
8N4Spkl4Ard3yBxjoiVyn5Vw3J5sLAXJuSqHNfJV3yUwP/Q/OiBo4PO9KD6WfZbSspa2cdBagI7w
nGAsM6OCUe6BBn4aqxYG1FgDwFC9aYIsy58poOyGReWQgN8gPHh4afp1mQO5OfK6C0JZILOb2Wn/
wReU90wiRx4WyCgKlmquSYW4avdlbLCRg7+dAo4XjA3COr6Etriej7iw+UlLRTlNmRXRAChvQFTZ
K932Ebq5wxXs/CDPAXLfT+nr+VAvLJOXHLrL1nqUlXvjKUH8y6DUBfdLTdmLAhIJkTQuFh8Ekfc9
K1why6F2OG+LXlzXDDF1+Q8e5m2/LgiWIgJUVsn124/sjdOWZ415haacp+ExYl/c1SmgTKvtGhDk
4Chx5UH2ELgb/OUCQRRJDdXqVKDDD5GVS5Y08FtALnwFqFIuiA/u5wEbq8pQ9xWCgqP03Lu/AU+a
g7LN/kv6+lpbgYhL39Wswwedd3JrqhMcsC1Mg665hKinbgSM+jQ84/xIn8B8muGJGqmMFwoJgwOG
J6XOzLbnV4+1t2zxKUCKxmiPl1HQutXDMSE4XqFtGAvIJ9Yd5dkdL8x04miMC7I4Lo25TFNCjWBa
z0vYREA+0YaaRXOmUj3X8wJ5+rNKj6cBwtwEDx63UO7zqODWOw2iM664+PaAgMcyRqpeG5M8Y/tW
fMYkTzFF2n67cgyPil73+Z9/CFCo44rgIDWMNJnt+LKUFolgE0Brv06n+xKiU75PsJEAd3VI2fvR
9kHbnCYLxTPwpYFzIYCz0kyykvO4Z7jHqzyvLwBYSA0mrK+JHcObJMVmFQuPbGVUC2IxEYGS5PDq
zOApVfi87Wk/HDLt8lxSHJLvYSvHgR1nHM01Myj96tFwSlsw9qXhZW2oMJXEHA99c26dsb2MIbKW
Y/jCIn0xgO4b/WqtBxtdSHD/dQAHE6BaEgofbB+N6sYdwIn8EyyajDxElpXihcAN5M4/kAUW6SHl
1CkYOrrtt68pHO9BZUZ+VBKQbHoeHWYpG5zDvhr+Ho67hYoh7qg/bMilA/Glb/sjLgKJkVvisyL2
H75bQydCzGRvKK6RmznWvBjmrFLjV1GmFSQlW4jn73ObcvkXCPSWBe34/amtyGVvqqNTLZ7P2+2O
POzsMMzUfhkh4eIOlGL4FERMzGyuUXlAqUGS32E8y4bQkwYIIYQHhE18NXcw23iIxZPsizPDdOhb
t9QY4AKqGWLZZplvxmT7xzGnnRvZd6sFoEWePMuw7di9VRCvAX/bTdCSXVUtE1TIaCNohoQ7T2Pl
rlnKtmapf4PhGM0y27yBVIpWUL1fiWpiSavHCYNkk3AatfruoIavXu6mdYQVrP6QFl5zRi8CzS5A
9dRA6xrsv0DczmFf4SFOApm5gjJg5Fuh5+pMn/rGcq2/1695uaEINs2GnbAeODA1iHj9wfd0KXNn
qjA9aJM3NoE32yyRsqxzmBni8TUOrKVDxjzgDE75LQhcBWrte4HH70PGkXT9p17Pha6OVVye+hwO
mMRHu/47V7Z+HilL7+HQMTR9OXD8rlvGtnTnzSXKW/dYD+aNXpomUG2tuy0iZR3apURbd8AKMPYp
v66DOOtGX+uazaZtY5mC+pEYak0IEDnSGdkya1WfqQZXZAtT9pc4pjrUCDquE697Tnnubu7Uk30z
770rLn1bwzY9LUpce/qp6/VouUDiMGh6SQw01rB69tcu+NCEf/8tebiDDLid3oy4nHm9QLTYtKyg
jzjVeyNg09czlQLc796ytxZJEAkl7BKqRYKJxkolBQXsjkFRv9loxNYpo5Jsd3cB5sxrL2wlWoZw
HdFLj3OAq518KYlqQMBUG/HKe56e9DGW+5ki5k+kLcEr2tKVU/o0hx8DjzHefHQAv+q5L8JiJgaS
oNqv8AGfl857W1hhRVMh4HscFgyit4HRXiSa3x97EPYiysoJU23sgjblxYScJyLElr1YHfz+/C//
7XuPI63VTZwh+FpLVQQmH+iF+0BDMpO9U67gk33Xu33fcTbbU321Y5ZxIyXIGiVujQcPFPVEtWZm
+eGdrWW/S67S9gAziN4kHmpyPgVWqWUL1DuIszaLa4NQE20YQRabCepFk6X2h9PveWRNKs/KXeyu
qKtXRz55eQv5T2WlcbPT2AZlO9S9q+0BTp/q4LPVxDwP8CBTyhUFR4fH0MsWY+XqSy7xuNKb68Yn
H1awblvwGtk/x9I1qFpJcCGIPcrD5Q81D/XH9fIQ1WYp0jPOIH8WRRH8GUwXOj7CvpgDlmhnL/6E
CYwvF2bSAlQhvANvZg63OGw2QDoNS7C4guc/azzVFr+aP8NOlGQmAh8ldOW52raV/0TbdbOEO0Tg
SxWJlJna3UJrruxDelzClT36a+H99WTF7ZxAngFaTd3oWYrUQZZgp8l5ZXlyegGMt998SyTJCVXV
ZYrUAXlmfkxHD1JUs7j6nKUi6Jdpop/tEIbiwyL6dJ9FtSXEhWCkcyJDlvlYbCNJYhKmf2KhU4VA
AxlOIGoqGj87jes5XoO7fmkPVMPSHQ9/N6ugwOOvZj1OXRHhQFQWV6zXmvNu/KWBkHckfKgTKn0I
5PGa+C0OzdbMp18WRrWNMwLX2/xwRm3ynj2yNHf4HyFOex1ypp8WlahBjNrBPfjWLEhJq4rAdGcO
uCDBHHoB7dlBetyQx60xj5V58hNEkYk2e4/jzE/OKO8F04aGAblmpig21UNpb/2ORwRqK7rYcxPI
VDmj8MMkn0UbO3wRdwHHp1HvJL9tsSxh37ROBkpt8bQnMyOy06aYtwG40yaFqYzdcL5+FWrkWO7U
J3fYBBUO6ynRQWYYCoojdoeqkYtOQMQN13X6Xrp2LqbNx6ao2HCWFQhJja1XKrPZFV6zO4n1Uzf9
GPnx48lF2mKHdtW53yw03msglXNayrE+TrU/S0d9QJpWtCwnP9JONIAAFf7BDvOem9Akoxv1KG07
aYcUM3aHt7sX3x+W/yc7fnj+AxWizcmPuQEDH5BkUMl8vASPgM4mPXXkTx7YhKtdCtptY/FYV97K
5lBrY0sua1sMqqgi4i7m6nZ7nznYcvs5SNcDU56DP1n7m/PLelhSVVUhoqcS2noGbdCv7b5p/9ib
NmXAzSH+BgePjZzKFhyWnvSfRrWEeCcnpLcrD6Ttxgz3aCJZ9BSpfvrQ82P7vN3ZmCZvPXlO4bxP
TeujkyAtRI1ZGWZyXDn0WF4g2aaMEYeo2uf+jBDXSXgEqDK844hCZrdhfJDM6QA14jRnCybejuet
iEK8ZO7qnruQehnmJ5KomfmSApIN11YTg1f8Ayc8xiTxno2nCKwyBzsu7k6fKnw/QjH9IigH85Qv
m15HEjVW2kste8DXjF1tsyiXOl6MtM9RJWOQOq+ebfRU0+qf658/bB2nxMTAG3y4oQDznLb+YSgB
Cyl+FaM6oUrJDw3k0IR8HAj33MaxfH3dcN5rkr9fwu0hRo9ijpyvhNIA6T26oe7CkufTav5s9b82
HDbNCdLkBqkUgpiz85ko6U9wqyA8Ri4cEMXPtkOrQoG8ihfilvWym1ZqSzLvVV8jaLTnK027900h
hPXxYB3j7XgH4hLJWK5Z70QLXUZEXl15+ZeRO4HDax9UcrxiC/eYKAS8DX8PqoFo07WmfG5UcbhS
OFm/d8TJ5mFYn1LQnUB7kn0SbwV3mwcGwbAUoBBhmMXR6/dEZEhLbOe2PBFWrwT1pmMTijH7g718
XtSN/PCEnym+G6n5b2nYptFHaAygSJtKbje9Ey7F32RvGCrlKMv4WSjexSOcaqIlCNk+pGAFNXfp
lBjX+mD5UdfFabAoLdFnI/1R93hGW/0A0X6zI9fzA+G3KNHoJp/dnc6sCP0AO8/aUbO88bG40Fjx
Bg9iUNn79hVvEkSCeuBw1JNRAc5OSxgco3iKhwSGEoEN/SS4fJWDe/qjtXdYDBfcyV0h7NU+gyQ5
b7Uf7qpBj22mDpoALw9VwiOqnOcgTxFfkT3NDV8tvovkjAdNFdmLn4taRE1t3c6cYRvP+6eyBjnX
mvcmdd7Q+o9rn3EF1j2MbWaFmbrzY+nngDimHmbVjpe/wUth0xCKsv8pCnHhpf1oOZR/eAvFhuSC
fdHnHidSJxasNVWa76Mot2md8h0K6RnQ+f1ty1PCRFURFqvooisHbW3ND/wRwZEgoinLXCfQiLPJ
A1BiuD5hX2k20GfcGhDBFwPdgwH2GLz8EmBJVNjv2hIGnwcnv/INjLbD9TUZcZcYLUCaxPYt0BUj
wp/50exXCwbM8eBT0+t1KbtY5/5fcOYs2aTmZZj2GBK0j8DYRw8NyEj4YfjoaKzpnI618U03ujNn
oR+BV9sKIfsIuG0rvGxDw7jO3yBbKEwmal/tbB8m72iFCNC4VFv1F3GTS0UWriQImba3h4rz0vQs
le1JaMSRv94DHfrUnickdJNCLRk/yNsb/sDwS6eqCs3C4i9o0NN3AGnh9oacx6iilqEC8TDyU3GI
hdemXYdlaiyKxVgNaVtn+4YpM8WZjdsJgHqs0etleWp5ZizSoiK+J/bK0wydvfua7DxTZli6iObF
GHsYIDSBQxZ3pMnSZdLzPSSlVwkWYJDrjbAV0rmUfEGtqZZmLgtUA4XJcI2lTvdjkAvbWqoEMR6Z
1NLi914QNifXBRlsgzl6QTaNBFdQVbfGr9uaN80kX+ASm1ty+slZ1geQVrMndZh8Dl+0km2FZv15
Y+T33/ekVUuR49N8dZev99hl5P1ouO430kgi9DH3z8P24VoNA6M17XB9Sr32BI+4tEe1W0QdcI6t
e5yQSfKD8FwgHQoNfeL+SsfEX99ffeEn4A/jVTuEUD/qCeFWB23rtyEmtUyp7/gkp0ffsy4JtC9j
qW60MgyhMMGLo6h1rHebtGZpuhJvNeWBtJ5LwlPZgAGKmFJTRz9fUaqQB0vmEc2vgfmOT/8IOjqs
5G/WHLDGWQMhDPPKuLyBCMYDealh4nQ36J+DD9ZLjLfSwjptkXavHvJiI/A3y2aaSqbnGZNwzcaK
bVfa1bSc9XaDDgIgcRILokD4ALhwXeG2J1M+FdBMhrunhLONZHDxWiro9j7WaIU//t4oMryMD8AB
xd6eehONz+UL186SekN84EmHf0NF1wyWtIFlvBJK92ZF4OcIAOUhrScXkAM7Q4QD6S7HenFAEEVq
lpQ6c7CBT0bIaPrLPLwEcrQPu9GACt2myIjJro6+hKkR51uF1T9NTTfpi3jdnaQW7YADFLewbFXr
DkPIEaEZtYqTVPNjc0nCtddWJ/zJ8/u4n4N98CP2zjLGDj+4rXcu421ybGGttpGs16H5LwXSFFbc
PJInisHtCyQHxcpnFIVHB/fCgq2HRlDlNw5XyXqux758WrTk2CvB/BCDUlubN2q8l1ttMWm6BMW0
Til2VMll74IDWK2JmyhlRPGAmP2IgPyNAMPYhtTltopEZ3peCkhOU9xogHHJbnjlZmhpFs+UtkPv
RtYVYhQg8+X1ObO2oTgaaZI4xyxgL8fPjnkVIlxYNOmEiSO0nQQic0qk8mQPDmGPjPUWGszI2Mme
1Q8sSZkg7PEndgI+BxZJhYGsyap/j0tsHFYGa36nK+3sivLbnTIqEIcFy+PUCTzMTB/h9QoXXKy/
fHwyOHo76cUaF4IDdmZUIXMMj1jQRxH9+cMmzgu1xIqoBFJNvNgUXoPBqstYl8jAlLbV0HGWXumc
2mVbNB9tuz+kwZn9fgrlDymBKeWj/YnWPkFYAXHHr4Tz5HyHzAVxQ2gkxsqhNAgTb0/LAj3Pf8Xv
E4oEtH2aZEDCMn0FkwkTyk8/7mVEdRcBnU03/O0vuVRUPdPREAocn6RZaGd9MgLv3yZPAK9leIj0
uvTZOaT/oMCzW7cTbu/NpxiLTgwV5/rYpRjKHIZmwVthQhLmVWj8P6Vq0bmu/2MuJ651ZCz467DR
u2f841yJTEVwihPW5SzP2gcZ9qR4ZcvO3exfy08SEj8rUV5vgV0VxekNFL6glDuIlrXpQCIDyh9r
rsXS+3lgU/Ol4UKSOQC4BbLr650Ot0NPRks8jpbJbH1ehVNF+amtnFT0YGG4JXMcu1e+3UomRLX5
LN6iWF5S+ls05PC3EvVYGn7vU5eZKHEwiklpT+Q6otcgWI0jhF5FfYnwxRR3LX4Ng51om1Vb6MwT
le050+FezlTsxDR9KGgwDB0Krk7c0KWq9hUSmni7rRUoQd3EQeUO1800p/yELbU5fWNcp/m8wEGW
ZAyGMoi3XfIOQi9MQOPMIYUzOxRNf9PQc1wAxR1pWInR/Xqsqx0ef3FlWcgw8niOpqEepI2tpbQD
d+CfFjPD7b3uC6kontznQGj49cxQtkwB6aAldOiDIsHDk6DeQ98YgdJddeLEaprI61Ppjj309anz
XBMraA30D3hnN3lpx8cR2EE5XWd5OYyABK1dCNMdiigvxsspk6qd3Fh7q7GTbdLwvdKCqbQiT6Go
TaZZM2LZZaMqHvadWvDfxlZqkz6c3q2IXRVpxS4HptSLhVo7uoAdqyPQldPtm8CWlt4UyJmPchYf
NZm1vkL99EnAAGxhioxe3MKt1Dz6YpMa1bHPriy0r8JJWBk5rUSsx3zpMBorAbswWcBXZfzjQ59I
zhaEAgHNlgc71j495ZYHLLXjPVfb5eUAFQbWYzrJAAEyFdsGP9l7SiaItRhODnq46KR/Bok+NUn5
GuYQEGU7EtiVpGbBAJhoUHuto2KsVZiwf1qeS5s1NOfUf3akdiAr91urQq4rA3/LJgnqCTFHJ/bl
ltvSfMsFeURWbHP21yWnpIS9TlunK/VyMJpFWbTEOJHp3zXmyGy3DJzIDmzUSaxM92M+zGG+c1uQ
X7xQXwDZxxByRScj9bfvQSD/WOGveIZ2sTJFvDX13T4SYtT2/pi/r2cioU4x8KEWDYnrI3WT4y7v
dDpZNy2KWwC/GA069DNzKHbdGXsOw0Do2zFq2dgPX84gMHtJCt/kYNGXYHnhmRg46+v+UbO0WbGU
8mBVp2qV1OlxL78s4sN3MRWUaplGtwa7sxPS4r11JwWB68kE04Kj2ePg8OxjKvu+lNG2h/azDq/q
0FbcPXVWh4cLc7zwDyrHjQtCtNOg8odVTcdRCy5UZj9ZpTD/jX26wt2CkERpSNqqYtEadyT7e48L
Uh8vcFti3MqJe+lIEJU/w9jQQ7PL0xMxkblWh03Z8Ye1vNJmdRLpzVPfgfU1IZRq8EIhmjZOzUbR
FwNKGHVzc7Q27DnqScscwalaN+JPG5WIhsdCmlzPIRE9UyF/ySVLmQwdXv/0d0jz4lVdt9/Dn8Cx
YvVgWr/Hf8gnhh8mZjn5FgUjeEO5rHF5nWSKmIDPPkvk7/sZIQxaww/iZpki4uIsBdYqA68EHJLq
jeAT5JCwJb5/OTTGqFmFpfyXyENeGXwIUi+v7yxG6zz7jEJf3cpTXiiC/n+V5ui/kSTjYkKq1sZV
guEZmS0+u/Lvm3jOiYOO1AWv1bIUBoh3Ve/9u/BbLY8xNImM1pTaW3biI9w2AVUJ6+LoliyXFUdw
QlwSmlMGSn8DoD4kJ+IUCWBM/c7LKevAq5SQGb1oKTKt9nNVHuEtruKDxYWVxHCw5aFwwWpvMxOX
Z6swx9qU3T3rOYo3p5D0plW1mKy8ifbB/GXNL19LXjsBxOeENT8HV6HxkJOxglsD48GAfgKs9a7N
TttyT27bMBgfSzP3QDd4FSg30sWIXeveoL2r22GFSg3IpwF6K7aMdhX7lWbpApFIfqq13C/9Gshf
Md6CjPgq6gGji7K7HaB3sKAKVYh1HSs45BwVqjdud5+gFWFzC1Rj8Ntn8mjq9hdJ8ShDZ1e37pLe
HWV2gqAm0Xx9+92d2OM528263bdP/AWOWb7fYkdAHTTLOXygYRCmvvEK2sO4WgbiqTvG+WnvmVyC
PYERLZvgwzhSsCy+OMo8pZFjyinGGzk1LUeZXhIg7zpuUgTjjEuskswlkMYbeVKj++k1KNe91sNo
/H1m67p6W4eu4ubK4lsr98+3R5I8EfzvvbedXEio+EZ1zDciZ1iZVfBhb2SkJtUQR5RPucDWyOdD
6Ngz9oGXZEzl3tgqn6YLuM6JEptaCZDIONh+rdtk1WDqmJv1ro86OGs2ZM/V1I5oyZkGiE5nqW7y
yNoqfI4Ojd/GXsIt/hANCCV5+FWzBIPGE9Y4c0HzBRwGZw7AzALcfczVZY5eVmtMrmu5L1osEn51
Uqz2c7uTN0O3k7BBwCSlS3VS90gegKeMJPwWTDlEiya5Juky67+z8U72TfGdNCBRM+mu/vPHM8X5
nAOvIV2XrS55SQn8PFZpowavzqCrZ8JmUiO1cX1hPn2RQF9d/WTZpFZ8z1zpjkZxIYLwlLneQxq4
E+j7n0+6NJ1AN6MwiNNETM38gVClqKDmrNBfs7SoxgGapWlRv4VU6Y9WkfC1uwLzEXUGa5QwqB0R
udtDEULEpvZ3KgSmIvtDE+tP4j3wg4EMZl9bB0KNVjzWpwuLH0bNJGlsrkEQyb6ItVNH8jndJted
fLVHdxAmONdvTcd3AWfU9adlU6wpMyds0icJwfVP7XdCqmSDWveKu5NkLlK59X+hOFJBpi/9mZYl
u0vPhoLYFI0Xh++Wym85WUidG0aSxgqMKhSkRhqmbhl6eTz8ow8I++ewdYzqsZRYtjGh3HpYVgFS
oDG1L3POHfuytu42kzKFr3pi5bWHXF74ZzNgB6XQS20VgSk883NfbmO2M4bBoUq2eaDI0db93r/f
XObADNDHyP7RmFcNLqaUnvVz+dfJy0RS6MR9CBWuw60frFiMwDu6SPEAQ+MgOsFr9Bna2DbwpEfy
aPAaDZ9IY95BbCA4WzHWJquhdXFYoymFtLQ10MLN3wnNoc7PUoQCiFxkATMvdf7+I/3UNujxec17
D7z4dfQPcr8zu7xM82OdxJZfqGovfZ7HbMR2KgRinngU1oem/uX+HJEyOIdP979tRoOnhglI8k8g
L0T6hGyKHh4a/FqaGPn8HzZRQmt7BSPtQc/SqJFn9xX+El4gWYi5TxOQfatgCgZ/mFZCgxTc+ok6
sc2OPrdL7BwNNaZgKGv5526qPBoIa0w6upymCb91Rgir7O9HSPlXcBM8sJONCdLcaUgBTANFtymA
jdhnfcQC0ZcrhKjEjU/tDnTAPZZaWVzKKbc8yfiXpNl+h6s6ACu0V3ZtYtACRln7L9BjtbeFiE/A
Di9htVZon6KANoi45EufVEhtn0FWG6QdwqHHCTDjvakybalG9q0YYEYNxjUyU5AwbiNGQLJ/S5fJ
VUU6n+Hdhea1nsJeJ4cvMEqUm+WDgrBU22vzrafUleljuapmTbUy39GNZ9JIXl5mtVaOeKOpwbjd
rT5dD8zU97evPnS2XvTG3wUG5+zZZ6/jfHAI1JUk+wwVS4j3B0MLDk3Uhjqr1zW9JWS3XF0ofxg/
a7uMfnbvDD4JWaX9Ab60OU5Hc8BLbApTVrAF0XIeXygVoTmRnW0AXlREZbaA5B0eHgpU19SKA0GB
FtYZDZNVfKSdHMtetqqddRRGSHdW3Jvove/6gTRthP2Ozt2UZ76sOtk+mUELulaUhhMJX5568x96
eNLbxv+Y5VObq/FLkKW8bsJosKSqmoOri57cG4rrbhkBMUvB9eh0qz96UCKfU3Gxi4ozonxwFcjL
qPu0+L/5SjW06vRWvl/CvUIO+Ll0tDKRFlQMz+VlUDWXRGvBs3XKsmIFlP4Uruf+kAs76SkIir1y
T2ogbf9eNjfPu6DAHsA5FOC3iD61ysMr4COD+ykqoAHi4MGbuSirthPIVEv/6hRKGEcnR2CT3Cjx
hVWkdqVw2wz3rbYa26xHOIWiQdkCgBkfu50ek9TAe6T1i96HgBW4OtYKwE/Qwi3aoT9y+g2SJRZA
vmJkW5Vfu5rChHBlO0wigubhwifU6QeGGz/f7rFczP8KTjyH2YQFh/tRy6wCfXlE6+xDJHd4rE2u
QflbCqDqNwvKY2DEz8YhHqU8+puC4RrIxNtqpNOnpElS2uQ2bm8XMV4LotRLaW9XlmbMb/btIA6o
BXyaDS34+yXQBPEkuODyYBAjPqWMU3h8y558CNVrbMFV719i2IEsqJHPCRXQ5moC5QQkaqCy233i
+I+k/OErUpzht7rheYGosbhFntDLUz9zPA4r/wpLeYgWwTiitwDh3tH/8Pf7Tzf8AYMNLHfOlDFR
Q6Vl9VdCgOooJG4yM3Mzx/AZevru2vS0gAKd9V0dAdGUKUNvWKRFqRavNv6R52BYxcLqu8dpDXmO
4olCDXGFHMCfo+YsCQB/vxxNpvCH7ZPRjKuWPiUmZBCaEU8QFHjo6MLSXg0VCQKdRh0Dhk/BQUbv
QkZWWZXApNlg0nco470Kkv/lvp/r9ElWIDWlb9I6Lm5chEKFgD2e4OUjbYWNzOmrQSPGHTQgxui6
26nTvgc4FiJc81UrEdl7wr+JsGXbdDeFBJm8l0SoVhw+SfMKOaMTE7eaGPGuKAqIEYOH+Yjf7773
u5F+rzGHwuFPJX3iHrvxMTkpLYfiZzALIw2Bj7jvU7qAQWr1U1a1fH/ujHTEw9ho7cGytTwqCTST
tdjy9jW6Y8FizhroWaF8Xqtki7TULsb8QjuRotW9B6DK0QRabztl2OV9pOn8bcGIfDLO/jLuvz05
eaqLhUvJaD5K61mrUEbAKeXdJvAuGixKQ7x3cMXz45BmXkTUXfXSoadOwQxt8Zcz8PjpNh+R3d13
3bJz43E6hqMmldGMkMFy/ukVLU2/7wdkia90iqcedPT549xAdNRq5Y8lqb0C+gQexsE3tYFFKp3K
qE1Kv/OqQmUJtWQnANSypfbtv+r4UAwqycPcXpHtTIN89Tg5hrtfVDHbq6d85Bd6Y7WepM8fFJbY
4H3LWWqQP2BSQiweUp2FeFfApvtnzmbbWEdIMNzcsOrfibsDrwfXnF/cwzR1ffzjzclHUWJzsprL
S+O/6/p3M0fyheEgscHTSAx7y/3P7GbOZh3lc1tdtspkFQHHNN2WjVQiCykYGbhtn37Tie9tMQoJ
P68syytGvpJTATQf27RRfXDiZcd2/Ib3NPxyZCgwy7BfYsUKdTCDTtH+GLAMfH04kB27od5e4Pg+
AFgUbylTL7Z8s7Z4uuj0cQWO5EF49eJ6yy9F1vL9ZM9DbxFLucB79UTjClvoa06vEZG6D8TDnRbV
rMtPWU0Vi1W1s489JNJx9RqGrOWTs6L7pMdp5BtXgJXjBm6t8utNLkfyWDhU1aKJW3+R58o6IGkq
xFEO0HeIAaj8xfo9+3NlnVP1/tdDONZvPEp2KgdMVgJgdkqfbICzC3v97Djk5V4X0nm3t2tDIItg
MQ9MjJd85aNnbRmA/VWpsXtaJa7G6Tzl0U5+5iy8jcz+ekckFTXGhow3lYPBI69VYLF2bl5VLTBn
FhJCiYqs6FjdTx378hkvMKvJEaluL7lniwLB6yNPjq8LfU+rp0/Af4pEQH/XXtwbfng3XicD3EN8
iTYh0fYNZNOtjRvRLz8Ds/7+2uYqlqYq4moc5Fzf6ctvvH3VhTZE662D7cuJeRag9G/yHP/+Tlw3
bfbNEwmU1yplm64vyVOAKJd1FF9uZz1rjQaZyt8zVcOREEC2OvF4VEnukGU02DfNO7di/mKoTg8L
Bv6DliAFt4KaiR/G9ATySt5CC7hgpC6QVzUpmASGTW5jF4kBhWyHNM/LHIoqThtP4TfxeAjVVKDL
nPGVW/n+qVxQ3fW6aTGgRe7twPMk5rYnDQGDjSzW5VHBQa4g4ukJwE7fUzEtk87NCyVpts+4Z2CA
WnJm/bsMD8aNTPPR5+ThlWyI/AvlrkznxxVWvsUyC2ibmCe0JzwOMXysy/dpaxtH3qMudmkuSnjX
Ov+toZC0EnNTJUMdcFV/69NKsSWJtr3x7YRtYqTphILPEwHaGc3d1gGUN1p+aP3tapfnfzGbTFrP
bGRH5aAzvj+WVNu5frxkhZq0PFkQNJh86RsKKCv+8Ek1WB97/ZJgmcQ2uegcI9qNTz5br0X7gNGj
j9KlxxPQqu0BVBM4mciYr0NvO0El+awJq3gElArp9x/6VhzNUvnKFsEdevKeYf1tub2+E4fTXnWd
sRCZPFvrl1zZuXRxNH21Hgmjmz3rBDMGxY68+cuzegchXjlUfPofSCrbYiclbG1xqMQ2X2k/hnqO
nsgkHRSei+WrfEIXfABOY3HObpcuzJp24Jk4Hm1pqC3GXDYeuQFpMozp3FiZrpgZkxhrMIarWkPQ
y6L7uRnQDQTvNxDfOe505Nn4adr7wFKn5vMFPTWQXmCoCbJe2/bxJhwC0GTINOk/tAbdhm5IkmJ6
ij8fITxJqOYQS6kON9BtNArNxlSklH0ERCJhWKzNyJesPfhZ1Ofv7GxR/9aj52anzb1RNpYOzfG9
//X1PM4FCFG62PEv3lOrzE/UhAgeGvtqWSKi3G/EalhSheTygIizLU/YpwJ07l2VBnp2NM/UKMsi
hnmSIRj0U+8X0vEf2xCUXmIvHri8CxK5QmoI2oXrsAZC4Ygzr9w6QumtQUn9yZBiDRUnu0H7phzl
URWGii/V9ifrLeYsQrmp4WtRPiAfGgGBo2CtPJo8NK+m0oCvCetA4THGRoZGO6627nOvu892QSlo
u2UDXGLBrOOD2G1ZBFcbZIK45IzO3nc1e2aRRUlmTPFLx3UQ2gGtYtRi7JnGkHhAjWrQx4vWfFjU
ZscXYimL8YvisowFEnExPJRbIGNlp9arNJFMD5qm8feufrklnNIPpsCcpeMDWXFcPqkkqO61bfLY
fApqlu98x6y+TSF6Ws5iWXjxV1QIvRabQbIwfyjXddXrTZKmuA7Z8pVNYLBBe2/btJdfrv8uT92k
ouVkFlpz+PeoodEXhIScpHTaZN9i5bkahpMirWxd9yK04ACMzVJLwOueiGlZfOniCz9ecfwK/DdL
z9qiSUy+fHwCmMJxROBkhhSVOhgMj768LoqeyjAYE+pFP0UO4+s8pHZtbnksy8Spv1x+kQ11o7Ag
nmfGYVbQHgywEbHYik2B40IT1KRQwUnNCMehBbAQWXgGIbJaqbXTUM/Z3OorciVaZfAn83i9rumB
Uqv+tr+X8PdcCV7dS3vSTrmaMSKc2UiKYBQvzK1Zyz6leDwN/6qXljDe0a+F6lk8NULoHqSlkVGr
MaDV81pusFdVPV3QJuTCCUNr7whM6Cpl8ROnM8Hol3cOyPKOGasbgl3D1oMpLZM9kYG+4VNg0HCc
GSIjH2h+ucG7oEyIrV9l9O57qFTtTsEXh9LxOz5C2NYMdBiS8yb+qfbbYq9RMt8uNFwZb1AeL7Ic
DeUw8fr2yZLgqbXjb0q236duzdQ5dfjHNR9Qstgj/NMggpgwD7ln/fXG+keMf1JrlpXOVlsr+iYq
l9ajC9xXRONjrxWOmONNLdRD7mem3LpDDz+4qshS5rP1rmsvwWnDTKrjIAXqKiiUF0cQlzVykRXP
NQ0EvSQsaf22IatBGiHw7m5rZ3DiThIOqDAuaW/7CS5sUxjknqkKnYIFrpyrD/GZM0BJtz9+3L3w
VCWLc9fYUxHej+U3xunxd7nsL6vtP/9ht2qIswAMbXqetIMpYYiy6C6x8oLDGwWd3bFLNXG+4G0a
38iMRX9r9lJW2ma8CCePduPw1EVyWnX8GvWwz1Mv0wxvbGZGc35frnt5DP7PJE0ZT2tDc/fRw1j5
6Az4efNugIeQobDUUFRu/YmZbcmJ/RYeilpanxm9yAOA6QeGreKobRav+9N+0uhRsUXRcRv+fE7D
yq5Zg0P8n/7ZlK0xrStisxS4HMrFcOFnFZaxWw1uBMHR0BuXTwwJR5xYix9Mdk1SvRFIPvNtVhUF
RUga37FnaWTXfULIt4wtmf9ZgegY9+j6SzFk9ltHK4SUcOKd5jICX9/Udixj+w7b7vRIMgrUj3fk
Fx4DdQRzQEBBHbozAgh0j7yhsOrqoq+XS7uubtqqIwsz0hofiMDtbgbxWcGZ2zp/5UlrvOKuwGOA
Ijg7LA0rGGWT3UtjyznFuYyndykJHAPU8ADpN0aZIaKFIfqLxzbgvU1gNukxvcHwCrviXf9gYp+a
M12llsQqLr22laCdJg6e/yoeE2/Xe7SWJQh91mXfE2ZopAJu1eFPeFVEbJ4AvqrRhGCMWtr6BGzC
gACPqb3UDUmsM04zVzwYVD2V+Ojga/h+l61TwNIh1YVM9Z9xNZh5IfJDcQrJuhBzWGLK6B7TsnnZ
9GJdDyjkjsagZBCjAyPr4VWeehBL0j1oRlHZ7Ioqt8TyLe87z1viSkl2d0lSQU7aXIc6qDuq0+mi
49/Kdqmw1DEhabszuo4vtX0CH4EgYBdf19fB02/2JBh+Iq+7fxANlIC9dPtF4CkeC8GPvbg2D2H1
v7a5ZejZ0ZaK5D9WDEADORh+RCFq0WFPYZjsFguOjL52qHcRMQy+N83t9r6DXLRCApuE92PrtjGD
fIK7eFSoprbOu15UV8umqNpWS/rc72AYeMkvNokdaPQYKA6S43dAf+T0/Hs5Viy46cIDEYfltlnA
Nr5RU5uIQSyfm9PpWySaEGH7r6otGzquFxWVsndenXi83cjMYZWhGD13Pl4N6orIxXXpjQDDMail
lR24BiHMGfm4Nt2jBIBBwTD5aGZ1ze/+Ga1mQW+h348euufu7MpjVuOdlSxmyx+eXXp43X9n0P4c
nsd/H9LdJFes2iBPzgr4n4QDmAsSZecMunDenPW2dCyMx4X9MWOpxiT7ibUPExrJN0U+Qpz3u7Yw
s+dWWGtvfhKmZJzjjkqSx6oUu/39+yq9E+GmyrEhliew/wl4/tuyMjrX+i2KYSx6OI6fJXVFVulI
djX0N+mvA6ISZoedDF3Hd1cBxtk8LkJbrs5gFpOeAc4u0olLb0QZXegbmbkqg2V6kT3a875w5vU6
Z+5bb6s56Iz1wkbZ8yFFeaQ0DshsUt6/25L2adOslvAaRanxtT6vcl+lGYykHg6rF1FdQrG/ziWi
omI2+4arGymcx1/1LQhHQJG0+ALc08SsM+/jb9U1MzPKFXmRysaIC3o1L/rCHlzhDWwCpTcB+AAp
btfHHDyPO5q4BzmNRHLV843KN2Do0XxJLSFHIu4YmrgAQ2y1/TH0Y7x1adVr0j3vpy5vfJtSdkGw
1YKVPqjehamGtYrzcy87ddCwqAHs0Ww5DzgGQCH3UgnjRCi53J02CNLZgLpGz0SOtoM6iJ4TX8ck
BSRTdJQ3RoYgOkzFcTyZaOcJyw/CrESsJUKCcfuL+heOFqsClIYrKn3wrPhYAXHkK4EI1jfdVCz2
bv9XFyiuYjJGunvAkF5c0nmGCKzBL5SWeq7H5wy8V251QYBoUd3UoKdlwZI2+p95jV53AEUgc87r
0JvW+YFkDdkhisMV4Gtt/MsBWby88pyDsP9XhGRr1FXsjscqJ6QehZzPOZVm6L/B69EU8YGTN3ww
XDsrrOR3gr9mq23pJFRzTTGznB57JKlIA2PsdyBZQYMlQqFftMhApNVVtWVOHHZQ78W0A1Ha8v4x
5E53o7QlqqoY/DyxrgWzWjpBXH3whPPJeLa4O2lBmTuT5QEx8/JQa2g1LPhBPwvsltsu/J9VOHZY
Z2mhTNa5/LW6IwMa+Q7SOijgOBf1zo3sYEJVdY6NhNxFTJOVanX+pd3F+Vh+X0CCCUUSOpdjOLGT
Rk1TaVtvfA4oePrR+2EH96cucAKLPQeq+XUPbp0x1EMeyX7CKFJpfZ30rjIIdVsOtNxhd96Zzunp
rStYyIaTcHzvIJgbdLYzl9M6rHbrl4eDKqZGTXfNetiXzg7gP8l9zdGq4gRuJMoCaq+x67u2UKQJ
cN3rOVYOKRKCwG7a4B07Mv7UQkD62WwdJCAWvgnS84bi9qS5lZ/3g9L8gwOg/gDVDkshydXLWvl0
+6mbbqsuRDdKzNb70WGYkwSd1LcIgHqhgLEWOvz3Ze31HP4j08nFIe267gUmWS391yGoZJ+gvKpc
YO5E96nbh7l4YYGnARrimQjQq3FfjRESfFThnJLQa8Os1nVCJmY5PZNt3tvykgzA2DFDKyfjFaxq
526Lno4PQZWiwmw6p2KiZNzhAGrZ+WQrOSEgeI4xOmPo45g4ccES7wmkcHj8cvn3/1xfx8/E/aHh
QD1fEqG3quTPvRoW+OjvI7QkaN8kql8JO7u1uz1keOG/fHDAlF2WtZEDJsyWCykTrxGlmlC5USy9
HJjPWyA5IvO3FeMJxO3Kd6UVAeAxYcgUKc3zD3mgxauzpsiyJKeY+Ku/ykMJIs6JWWaqmXcDoqkV
S1rBeDahiswK76leqqL7ESS+HxxsVR6m9XDhI6FXDhSMdjDLLElA4TVRQPgSrnN+a9ijIX6XQ8VI
QueWiQzEOi2ULVC136DlqA5WzRC07HKDVv8h1uSGbLg238eMB2K44xRB712jIPCXqXV4PlnotRRF
Jiy0H5j7iN1+k/+U6aoznxfdZPw8XOLMbA2dySV2fhJwUFkR4J2l2ENOqPliVuajdhsYjgiDpyTO
yzI+IIP5Mqf8Ct7YHSoZaUdNI9gXYt/NxvfkuVwyRf/Sx+2TEl9ngiEuuJvh4oRwR6KwONthSWjY
C5LWnghjb0jM9eDVWTdhUqMyKwFdeRYZHptf7pUB3kM79xJ/zVdCXVVpcSKF2noHx9oN+sIHP5YA
9NChOYnMsajmWyk5aJA9H5aVWQOere3cGKGHX7dhIbwjuhbkql1eDhHHuIHvifu+RnYJEuQuiz5F
9eKQRKi5QiGAgziksHkvrzhRbHec7Uo1k8rR0OGmfE1Apmc4cuXHwFRx/VKo/hOr8w1VpeYAzUQj
tb4oOTkwekOXR8gaF5oUR75YCu52xx4ylNQ3Un1nOB2DCYKysMggOPdVWbhEUn0kV20L74fMFxVp
qKFgLJDCIiZLgXtARSe/EpXgBnac+cM32LjmZZ1fI953K4R0VaMZ3wDLv/3oQ+GeAFWs1OzajY/o
86XfqN0pM0OTIWmar2XqTM850/WE9YmyhBK0OIPau1+QnvLOstIS/0FIZITrAagIsP7xxe+TS03+
3tBdXlTPenaPFH6SPqFgsicQQPhLZ+O0s7W7CGTUoDnvQK8pjs76g25VwKO55EQpCTrW8arHCgBM
tkX9R58HIuzGb04thPE8yZglSfbKRNKOA2U5VHOY4yZnvpJMZOkA4BWEmD/d0q/nhlgBgBzokFUy
L/bw4zTufQQcrvY/OAJJwGqZEy0HRdFMUFgzbJlvxFIZ2YzJfY827dC7O6rA8uVCZf7VpeKJB6Pt
Z4lS7vz1bdw+02B4OJAuWM4qg7G8N6CY2SLbgzAiDVBMJ9qOS3GFvziouY3+K6PK9BEL1j2dLH3I
9ywCKxekEiW/nkIsFGNIPe6Ams05UNh0BDfJ4D9zu367Hbq8JJBLf/F3ZI08rYxj5Y+OBeFh6inH
vPMtRSUzeXhd9pvJPSwCPto543VOmITRYzCTt6pRRJ0R0ST2ec0oxl9EQxlzQaIIqOgNGIB0CoYz
GD8klowNhLVqp2K24Ct+wzjjQzEPGMxkwJM7jsdmJ/Gm8DC7N/oHTViRNXD8mdgL/tls4Ek8wTMB
MaI+NggjOiNIDLZWyAz2n2VZN45WD83PYhtNqpBgORv5f333jc4td92utF4ePiwt0xq/WsJOEvHx
3geAbw6EX5sZUxf0Hs/Yxi9dtswV1JdhLWjPxoF2eKIzeETpNvwCKLSwDJ2p3b9xOtcuv6BqpurW
5hlo0Ut1X/PNAYEQ0s6yL6qtmd2cnL9A1jUinAfy+pm64BrFeujdjYS6m+obdlvaMIea0ZCgQHUD
eV8kg4rYSf6k9kBbMp6TyhQRry6nyUCiOA7h1gLKfIyKYUqNN8aROibtcLe6bP2AfOBS4CG9L0J+
GTGZY/nUAUCJ/zouYL2zmYRxdOE44WuqXgZwf6FfwPEmcuornhzeT/xU2umktH55IkmjT4m0YKEA
hdjXKhnlrQKXQJ5/SFMxrjbqbK0F1xKO3hEto2nTQsM3dEbR8GkyKyvAnUdvud9rOLYPL4y7MJTa
f5DBpfiRM0k+2xECfDTPe3RfSqGQYGbcz8YFdbZBeIn6xPrjoKoKyxSKvVz4Lh97g7qwVaOd0FFX
PF9B9H8cPSCblUJZRp6OqbYcTtiRQZIP3C8KwTl2MYjW7krgnNuaODuPy/kRJRzjT8/KhruqUijM
jZ/uRJWRqU+Dp8tyRFq62uOXv0ZU1HuEQ0IxD/bgNOWPTkPMivnshdRiqpAQatxTAxsHOE1jq8n6
stOcNt8exb8kWnQhcw7PzcyVGlOzod+kzL109fmlaEJ7lLEdBcybl7/j9jThcAjicQM0o9Ybnnch
WG3TDoWFeGIGhQAs5y8B/b95ba9ojATPyi6WlgjtKFNZnqeos/nYOgRBLze7WAF2VEJNtIqDjYRJ
8MYMLp6nvtG/7StDtqdAtZ4eGt8neWhb4Yq3bIpfXj7MtY04eZP5QN6mDFsIY/yL7smABoIcq9LW
0VOicBV+bqSh8VMYOq5ZGKD2hzsaD/NkgJXsI1eSMUm6pYhN1ruQICJonEpj/pjQKGIEN61MigDx
UQM5f2vt3HLcl6/VoJa2gC+HcuNZm0FlJZkB4DTe4+sfbnDoPJPytGSsGUz1mMkgHKNRfQ5WsPMx
iUWn6vAbPl0TmgzRPTkej9K+d6nmiH5Wt+uroNVdo+dVSZoy8KhTXelAt8IycUYDhBKy+nm4PA5Q
W1D7sQVFTW/wKVRV6HhDKccFe7gyTskOzexUqDbdwOkVvL9NorQ2VwC/NPvCMA4tlINFCB6fFQI2
TZRmk6hqDdI0v6WHkKyrcd8XjFYfpYkGxNL8uP2lCVaLA4WMoBH9wkMqxmTeOLRSKyQvafnRxUVA
QoPdFAzMga3i3euC1hYIkioYGr8PhfMf7bM63mSlCYmO2ogBFnZtNdLaDdhr4xCsAFX3BhD4lzQa
O3GC48pLktlWGaEzS/QrqFqZUlNgPS7ii+fYXHdu4meOWrvddDw6XRyocREC/g8Oe4fJs7SPHX05
miHkrGu5or/BHuBxq0nrPfAxMPFBATGpPtichPmBoskq6EGPIV103DO3jnGWAyhPemp+ZJ7/eh7r
1HznZ7zGuSlXjGDotYBgqzEKKLT1iqKVXQz0obt3+fBFm+S2lkAXJghaZMZe+T0COEI1JEc1561f
YTVgHjfBteYp6oVUZsQivFy+gDb10Bgb2VoxWE4fdZZNg1s2X9JKdvusdrdwa0z+G2iDC2GFWNf0
yTIu2yBhiFNxCvYJHHj5u0gxMlW+DJrmnU3yQg1GdBkrK/jMz4IQ3oOVJn4YacQflKS4hMM6TzFR
uQ/lPNdtze+Ow+jxxU+mpCP68iqRSBWjm5u8vXJ1u2zmm8CtDovsIbjbVAA8N22idtXSXI/iH7Nd
Y1HPDEGZx3VucMUqd/EiDMB+eX3ZS2qIjI3n3G8NZdxdjXqqQpptr70/uiwmeOB49n308SgbQDOU
J08yodsiVyoZu5qg4ok416BKBG5b7s9MZ2Dmjx+bmBbHYooQ7rApQaJkZ82pJT0xST6lFuV9syxB
f1DFgFeIuucVkSK+eclGA/DaB0gDbcWtPOnf0anGgiPJRxAxmpQuMh6uU+0o4I5dUL+8G0wgcwct
MuOqgl0awSlir0Jx7W1hXNt099W+YXzvBS+Y1LGdkSaVh+OoCgY6WY3h60LSpMh2S8wEHRZhpnOe
amvc4b5klP76kM6UxAUXrzRJN/hx40IPvcj7k63Z2UFwY/nNzTSVVE4HsAvVqwqoYGZ/oGeHwlft
amIpDqb5TB8lV4LZjAB2LU2me5XXTA/aKZgU4jgnEcPCMAmKZmFO7XRtFexdXfPBeLLJd6bnI1HX
yj7N9eq1WXheLd1kzOXUhZ1V84YSfw79cPZp0eCrvVjFEQbPkIuJDySZteCMB1YGDAVsNogR5IIV
Z+jxRxqsqagPGZYuKTdHf/d+BzttlaGms6knqThI9rA5pEjjsOq0+W0ALDe/Dp8uOBE8G+crgA0r
XQNZ+23cQZoWkQ/70vRqe5STHLCBn7TWmd7bjR/WyBPCEyw/CSDr6Qki4BihB9vo06EWcWWVY4zZ
dpY8FWBsL4gQXRs7RVOFGA8uwkrZiiR48mcjADQnWSRkl64B0YGqTVIoVxJtM7dbqbjdbyktgAt3
3sNMvd2ugMFjszkagU3e43hEJMzUTCS4WlDdVnJNS756GGAeU3zRWDfaXIKgKPDls0YBxI90LVcn
AYAFSLwvjhmodftIx18/UUeyT4SsI0bOLcCOpiKHIuNcplrI9RN3SpUNrCY4TFrZNE0DFi+ZsBVG
NpYd0+aFlyM6J0FMl2Kxy4nHKQQ5JQaAf4ZBFNZUDZDcXnCYQ4FeO21IQljbhDymfHMMffXS7YRo
Jmw1i3FmUPpL9qmAUpoUFarfpxPl36/LLET3kUBPEd/hWh56zVvNfJ1t/i9ZOdabHdAuQUY6l5ZN
M/FfxsMoSFzi5V5r6cej3Dpf1dud5sMSgZVpLDvN8e25AYruRS0/KOn3rW87CJzicXw0MVL/UDJa
r3GCA95QEyDpvof6yrXlltwIh+iuRXJlwcbAXL8gdUAkq+wd5c6j1vSYysXZ5vkTCzz8GSDn72gx
LJuAtxICfmM6guO+iBRj+zQ2ReX9ijdIYmCBjUHPRnJxM8K25aFpEcg2hY7e9x9pkhAbH+biAsf6
ZvNkzhdAwKTKN/dizuR9gPqEzH7b/0GnZzrPVSuuBMQeDw4VxUrG89Eqhk+hdGggJGHYjReg428P
481h2bfSxuwG8VN5bkhCW4cjNCU0+7QoKfeMb31AIjQvowjM28c4ODm4FIXdM5ggAwbOZjtXZORK
rPRT9K8n0KUx31vHHECRawHf1kWOsDeEFkPISUXPs20f30kV1Df/2N+CCbdREYot1T96vFZqzpPp
1I1wwtzX3/rgQmJ9r2WneOOq+Js8G2pRFvgbctPuraYw6F8pjjkHpj8Dtm4/nMurXWyc+BUW0fO7
S0CpSHNMO/lILoq8lv4npBN3p9yuudBO5FdM9PKYdblydy7Tlro3WD1zXScQEOAKbNZdD7ZBtgh3
MMJZonABXwVAN8SscHDuEX0LTEfKuB820evFvPJ8oWDGjo9256uiFwIBtYD+XAK2/VFfZ2+c0G61
Nl5e7xyxZqm9J47kQwZS+bYbNVX9yeRNo76OX9f0O7hyP0D5XLbapDXWRhALCZ9ldOXTfMaOpVyv
pP78LkqbRqXqsinxSRoSiWsAeXILQvtUsWUGxACiN3WPfS1dM6cC+zwLz5kQdms0FjfQnv5hFFa8
1uXZPspFXw+6pHl6X1P8KHzT4WayJgrok9JJrUX33qSVuCOeiErE1DxwQ6i4jDSKjtDZkpQNvnKa
t4/hJXDyQ4cdg06GDF9PKU2oeEudpjEtHcKOObDdm3BiV2DQOFDsSIM68EaGrIYJD0StpHuPtLco
cngMdxxLS/6um0yxlxcJ3at+riuZLsSfF/DiS/SLv/EPdy5T2MmnqUIOAW/ojXfM06bab1UP3+qz
2t/wpZf+Ab6Zi17wvKj0CXFyneoeWKt265NTJD5sMUYtuuU8FABVuFqTrrv6cDiZ+aLTc/5StVp2
RRRp4uFY5c4Ma8nRKDjpMg/CYaaswoE2HYBpvgpTOK+Zu2VNFBOo9cC6vsLHvvGO6/IO38lCjIyH
4ImgSdVNTTALhbz50HjlAVfyO8mSYPnFgQj2Xb3ZlOrQdzFG764Fd7PyW6vh4KD0CtvVswR/R2EK
+5MkV2yhXAORLAeKWLNUg2mQUZnIO+rHOnwLJkuKhDvn7cwmcoEtjwzxnDxv2IwnzPY1zzOvLA4J
BYfYNiDIDq0q8L8x6MRYF2ilnZraY7phy6Hjob6FiikbgFpYy2DevbG7Z0Fd7Bn6H0ZCtoh03maN
oaOaVHwp4DhYKIB9fCG784iGtPHWYBRKzCYvC3d3kxMgcUW8xgsz9v77ZlKOBfOvUzdYuzrYP/+X
r1I8rV0fsGXl2wBC4eGeP18ALNxb8h5HfCckkMp6hDU8ujZQ2ja14YO2Daz+dp3MtTFEEQEXNuo9
WnOKMxCB0AnmkwAKTsCy32IusUFjxxJULKDjd6duIeTOPAAQdtZrBNL1NJVYCxPFiw8uGwPtiEL9
Oz6kNKXv2QQwIhiRqn1+wZPt4fSHsZDAm+3n56PtMU58n/31NyvPrn76aO8Khb2cUBZDolWaEQcN
N1SFupxTuh6xBBCd1T4FLos01/VyQNmCKhep0yb3T4l8dJKoCdVRjRQyj8tqdXeeeAXHP2osCqe8
GD6g9zwUMwAyZ8gZnjraG01IJz5wyp2XgZEhA2vL76w2AN2IPs+tywZEFql5Nqwr7x2WoAz7wciM
2t/kQ+MdO6bJeo+1a3UEe2uKLDpFevP9mV585/K8vYKOwnCR/hLI5xkOEmw7p+f8uPdw8SlkvIzT
6dhrOgnNAvmwdGb6J3/Gpjf4Ja4nbzJvKtScbT25brYmTLQifmQQIsmM0q3rqJpEk4W/GEHE8Uz5
y57KwUMLyiSHAqLqHjkFH+Qnccz6YAMLHMStDqarmLuZwBKR5Y6o0+BcZ/tGB1W7a0XGS0jNMN4K
5hBM8rJJvQs82l4KII/bqVzvlEDS5pu599+uF7N+rSs26kRWJMfHyBPP7ehV0Gjlyc2xYLF1rgHA
Llx727pAwIiY5Q0wqkFySVgplE/EswAtgzQt4qChF2nhnVO4VpBIBVoMycOPqc+sQ3ET6kDqZ3SH
RAXe9peZe/L8KhZ4smQnM9CmJ85Ey2oZUxrAvSKa9kdY2Rl4UEerAz6pbjH8rRupw/eM+LoezM4t
RZX6X9XgeGGLzw+WTQFe/DN7nEDuw8lycgs7/Gr8j1O/VGcowNbtxLzVt8eEQf3gIrbaVLod0ykG
PFdxjdccpuiFlgtGS3XUCv9Q+btWXkPozd47iFo0wzzr8Erb7V+F8lP0FutOszru9C1dA1Dm/lOC
bNi6KImpMW6KbSUUJ/AqVu5vSzoBliZH75zmiBIVBge6vTGcKD5yltrzouctbjvJPOKYYrW2/4GW
8R5SHnxc3+xcFR8BBoSkPMOKoHChYCTSBCMG02/m0bQ0VQSnG6xnez27Do+Kok5/LVmw0IKV0lxy
am4mPxJxXw==
`protect end_protected

